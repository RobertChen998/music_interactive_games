module color_palette(output reg [23:0] color_map [0:15]);
    initial begin
        color_map[0] = 24'h040404;
        color_map[1] = 24'hf8f8f8;
        color_map[2] = 24'h787878;
        color_map[3] = 24'hd3d3d3;
        color_map[4] = 24'h3c3c3c;
        color_map[5] = 24'h8e8e8e;
        color_map[6] = 24'h272727;
        color_map[7] = 24'h000000;
        color_map[8] = 24'haeaeae;
        color_map[9] = 24'h535353;
        color_map[10] = 24'h696969;
        color_map[11] = 24'he9e9e9;
        color_map[12] = 24'hbfbfbf;
        color_map[13] = 24'hfefefe;
        color_map[14] = 24'h161616;
        color_map[15] = 24'ha1a1a1;
    end
endmodule

module image_data_original(output reg [3:0] pixel_data [0:59][0:59]);
    initial begin
        pixel_data[0][0] = 4'b0111; // x=0, y=0
        pixel_data[0][1] = 4'b0111; // x=1, y=0
        pixel_data[0][2] = 4'b0111; // x=2, y=0
        pixel_data[0][3] = 4'b0111; // x=3, y=0
        pixel_data[0][4] = 4'b0111; // x=4, y=0
        pixel_data[0][5] = 4'b0111; // x=5, y=0
        pixel_data[0][6] = 4'b0111; // x=6, y=0
        pixel_data[0][7] = 4'b0111; // x=7, y=0
        pixel_data[0][8] = 4'b0111; // x=8, y=0
        pixel_data[0][9] = 4'b0111; // x=9, y=0
        pixel_data[0][10] = 4'b0111; // x=10, y=0
        pixel_data[0][11] = 4'b0111; // x=11, y=0
        pixel_data[0][12] = 4'b0111; // x=12, y=0
        pixel_data[0][13] = 4'b0111; // x=13, y=0
        pixel_data[0][14] = 4'b0111; // x=14, y=0
        pixel_data[0][15] = 4'b0111; // x=15, y=0
        pixel_data[0][16] = 4'b0111; // x=16, y=0
        pixel_data[0][17] = 4'b0111; // x=17, y=0
        pixel_data[0][18] = 4'b0111; // x=18, y=0
        pixel_data[0][19] = 4'b0111; // x=19, y=0
        pixel_data[0][20] = 4'b0111; // x=20, y=0
        pixel_data[0][21] = 4'b0111; // x=21, y=0
        pixel_data[0][22] = 4'b0111; // x=22, y=0
        pixel_data[0][23] = 4'b0111; // x=23, y=0
        pixel_data[0][24] = 4'b0111; // x=24, y=0
        pixel_data[0][25] = 4'b0111; // x=25, y=0
        pixel_data[0][26] = 4'b0111; // x=26, y=0
        pixel_data[0][27] = 4'b0111; // x=27, y=0
        pixel_data[0][28] = 4'b0111; // x=28, y=0
        pixel_data[0][29] = 4'b0111; // x=29, y=0
        pixel_data[0][30] = 4'b0111; // x=30, y=0
        pixel_data[0][31] = 4'b0111; // x=31, y=0
        pixel_data[0][32] = 4'b0111; // x=32, y=0
        pixel_data[0][33] = 4'b0111; // x=33, y=0
        pixel_data[0][34] = 4'b0111; // x=34, y=0
        pixel_data[0][35] = 4'b0111; // x=35, y=0
        pixel_data[0][36] = 4'b0111; // x=36, y=0
        pixel_data[0][37] = 4'b0111; // x=37, y=0
        pixel_data[0][38] = 4'b0111; // x=38, y=0
        pixel_data[0][39] = 4'b0111; // x=39, y=0
        pixel_data[0][40] = 4'b0111; // x=40, y=0
        pixel_data[0][41] = 4'b0111; // x=41, y=0
        pixel_data[0][42] = 4'b0111; // x=42, y=0
        pixel_data[0][43] = 4'b0111; // x=43, y=0
        pixel_data[0][44] = 4'b0111; // x=44, y=0
        pixel_data[0][45] = 4'b0111; // x=45, y=0
        pixel_data[0][46] = 4'b0111; // x=46, y=0
        pixel_data[0][47] = 4'b0111; // x=47, y=0
        pixel_data[0][48] = 4'b0111; // x=48, y=0
        pixel_data[0][49] = 4'b0111; // x=49, y=0
        pixel_data[0][50] = 4'b0111; // x=50, y=0
        pixel_data[0][51] = 4'b0111; // x=51, y=0
        pixel_data[0][52] = 4'b0111; // x=52, y=0
        pixel_data[0][53] = 4'b0111; // x=53, y=0
        pixel_data[0][54] = 4'b0111; // x=54, y=0
        pixel_data[0][55] = 4'b0111; // x=55, y=0
        pixel_data[0][56] = 4'b0111; // x=56, y=0
        pixel_data[0][57] = 4'b0111; // x=57, y=0
        pixel_data[0][58] = 4'b0111; // x=58, y=0
        pixel_data[0][59] = 4'b0111; // x=59, y=0
        pixel_data[0][60] = 4'b0111; // x=60, y=0
        pixel_data[0][61] = 4'b0111; // x=61, y=0
        pixel_data[0][62] = 4'b0111; // x=62, y=0
        pixel_data[0][63] = 4'b0111; // x=63, y=0
        pixel_data[0][64] = 4'b0111; // x=64, y=0
        pixel_data[0][65] = 4'b0111; // x=65, y=0
        pixel_data[0][66] = 4'b0111; // x=66, y=0
        pixel_data[0][67] = 4'b0111; // x=67, y=0
        pixel_data[0][68] = 4'b0111; // x=68, y=0
        pixel_data[0][69] = 4'b0111; // x=69, y=0
        pixel_data[0][70] = 4'b0111; // x=70, y=0
        pixel_data[0][71] = 4'b0111; // x=71, y=0
        pixel_data[0][72] = 4'b0111; // x=72, y=0
        pixel_data[0][73] = 4'b0111; // x=73, y=0
        pixel_data[0][74] = 4'b0111; // x=74, y=0
        pixel_data[0][75] = 4'b0111; // x=75, y=0
        pixel_data[0][76] = 4'b0111; // x=76, y=0
        pixel_data[0][77] = 4'b0111; // x=77, y=0
        pixel_data[0][78] = 4'b0111; // x=78, y=0
        pixel_data[0][79] = 4'b0111; // x=79, y=0
        pixel_data[0][80] = 4'b0111; // x=80, y=0
        pixel_data[0][81] = 4'b0111; // x=81, y=0
        pixel_data[0][82] = 4'b0111; // x=82, y=0
        pixel_data[0][83] = 4'b0111; // x=83, y=0
        pixel_data[0][84] = 4'b0111; // x=84, y=0
        pixel_data[0][85] = 4'b0111; // x=85, y=0
        pixel_data[0][86] = 4'b0111; // x=86, y=0
        pixel_data[0][87] = 4'b0111; // x=87, y=0
        pixel_data[0][88] = 4'b0111; // x=88, y=0
        pixel_data[0][89] = 4'b0111; // x=89, y=0
        pixel_data[0][90] = 4'b0111; // x=90, y=0
        pixel_data[0][91] = 4'b0111; // x=91, y=0
        pixel_data[0][92] = 4'b0111; // x=92, y=0
        pixel_data[0][93] = 4'b0111; // x=93, y=0
        pixel_data[0][94] = 4'b0111; // x=94, y=0
        pixel_data[0][95] = 4'b0111; // x=95, y=0
        pixel_data[0][96] = 4'b0111; // x=96, y=0
        pixel_data[0][97] = 4'b0111; // x=97, y=0
        pixel_data[0][98] = 4'b0111; // x=98, y=0
        pixel_data[0][99] = 4'b0111; // x=99, y=0
        pixel_data[0][100] = 4'b0111; // x=100, y=0
        pixel_data[0][101] = 4'b0111; // x=101, y=0
        pixel_data[0][102] = 4'b0111; // x=102, y=0
        pixel_data[0][103] = 4'b0111; // x=103, y=0
        pixel_data[0][104] = 4'b0111; // x=104, y=0
        pixel_data[0][105] = 4'b0111; // x=105, y=0
        pixel_data[0][106] = 4'b0111; // x=106, y=0
        pixel_data[0][107] = 4'b0111; // x=107, y=0
        pixel_data[0][108] = 4'b0111; // x=108, y=0
        pixel_data[0][109] = 4'b0111; // x=109, y=0
        pixel_data[0][110] = 4'b0111; // x=110, y=0
        pixel_data[0][111] = 4'b0111; // x=111, y=0
        pixel_data[0][112] = 4'b0111; // x=112, y=0
        pixel_data[0][113] = 4'b0111; // x=113, y=0
        pixel_data[0][114] = 4'b0111; // x=114, y=0
        pixel_data[0][115] = 4'b0111; // x=115, y=0
        pixel_data[0][116] = 4'b0111; // x=116, y=0
        pixel_data[0][117] = 4'b0111; // x=117, y=0
        pixel_data[0][118] = 4'b0111; // x=118, y=0
        pixel_data[0][119] = 4'b0111; // x=119, y=0
        pixel_data[0][120] = 4'b0111; // x=120, y=0
        pixel_data[0][121] = 4'b0111; // x=121, y=0
        pixel_data[0][122] = 4'b0111; // x=122, y=0
        pixel_data[0][123] = 4'b0111; // x=123, y=0
        pixel_data[0][124] = 4'b0111; // x=124, y=0
        pixel_data[0][125] = 4'b0111; // x=125, y=0
        pixel_data[0][126] = 4'b0111; // x=126, y=0
        pixel_data[0][127] = 4'b0111; // x=127, y=0
        pixel_data[0][128] = 4'b0111; // x=128, y=0
        pixel_data[0][129] = 4'b0111; // x=129, y=0
        pixel_data[0][130] = 4'b0111; // x=130, y=0
        pixel_data[0][131] = 4'b0111; // x=131, y=0
        pixel_data[0][132] = 4'b0111; // x=132, y=0
        pixel_data[0][133] = 4'b0111; // x=133, y=0
        pixel_data[0][134] = 4'b0111; // x=134, y=0
        pixel_data[0][135] = 4'b0111; // x=135, y=0
        pixel_data[0][136] = 4'b0111; // x=136, y=0
        pixel_data[0][137] = 4'b0111; // x=137, y=0
        pixel_data[0][138] = 4'b0111; // x=138, y=0
        pixel_data[0][139] = 4'b0111; // x=139, y=0
        pixel_data[0][140] = 4'b0111; // x=140, y=0
        pixel_data[0][141] = 4'b0111; // x=141, y=0
        pixel_data[0][142] = 4'b0111; // x=142, y=0
        pixel_data[0][143] = 4'b0111; // x=143, y=0
        pixel_data[0][144] = 4'b0111; // x=144, y=0
        pixel_data[0][145] = 4'b0111; // x=145, y=0
        pixel_data[0][146] = 4'b0111; // x=146, y=0
        pixel_data[0][147] = 4'b0111; // x=147, y=0
        pixel_data[0][148] = 4'b0111; // x=148, y=0
        pixel_data[0][149] = 4'b0111; // x=149, y=0
        pixel_data[0][150] = 4'b0111; // x=150, y=0
        pixel_data[0][151] = 4'b0111; // x=151, y=0
        pixel_data[0][152] = 4'b0111; // x=152, y=0
        pixel_data[0][153] = 4'b0111; // x=153, y=0
        pixel_data[0][154] = 4'b0111; // x=154, y=0
        pixel_data[0][155] = 4'b0111; // x=155, y=0
        pixel_data[0][156] = 4'b0111; // x=156, y=0
        pixel_data[0][157] = 4'b0111; // x=157, y=0
        pixel_data[0][158] = 4'b0111; // x=158, y=0
        pixel_data[0][159] = 4'b0111; // x=159, y=0
        pixel_data[0][160] = 4'b0111; // x=160, y=0
        pixel_data[0][161] = 4'b0111; // x=161, y=0
        pixel_data[0][162] = 4'b0111; // x=162, y=0
        pixel_data[0][163] = 4'b0111; // x=163, y=0
        pixel_data[0][164] = 4'b0111; // x=164, y=0
        pixel_data[0][165] = 4'b0111; // x=165, y=0
        pixel_data[0][166] = 4'b0111; // x=166, y=0
        pixel_data[0][167] = 4'b0111; // x=167, y=0
        pixel_data[0][168] = 4'b0111; // x=168, y=0
        pixel_data[0][169] = 4'b0111; // x=169, y=0
        pixel_data[0][170] = 4'b0111; // x=170, y=0
        pixel_data[0][171] = 4'b0111; // x=171, y=0
        pixel_data[0][172] = 4'b0111; // x=172, y=0
        pixel_data[0][173] = 4'b0111; // x=173, y=0
        pixel_data[0][174] = 4'b0111; // x=174, y=0
        pixel_data[0][175] = 4'b0111; // x=175, y=0
        pixel_data[0][176] = 4'b0111; // x=176, y=0
        pixel_data[0][177] = 4'b0111; // x=177, y=0
        pixel_data[0][178] = 4'b0111; // x=178, y=0
        pixel_data[0][179] = 4'b0111; // x=179, y=0
        pixel_data[1][0] = 4'b0111; // x=0, y=1
        pixel_data[1][1] = 4'b0111; // x=1, y=1
        pixel_data[1][2] = 4'b0111; // x=2, y=1
        pixel_data[1][3] = 4'b0111; // x=3, y=1
        pixel_data[1][4] = 4'b0111; // x=4, y=1
        pixel_data[1][5] = 4'b0111; // x=5, y=1
        pixel_data[1][6] = 4'b0111; // x=6, y=1
        pixel_data[1][7] = 4'b0111; // x=7, y=1
        pixel_data[1][8] = 4'b0111; // x=8, y=1
        pixel_data[1][9] = 4'b0111; // x=9, y=1
        pixel_data[1][10] = 4'b0111; // x=10, y=1
        pixel_data[1][11] = 4'b0111; // x=11, y=1
        pixel_data[1][12] = 4'b0111; // x=12, y=1
        pixel_data[1][13] = 4'b0111; // x=13, y=1
        pixel_data[1][14] = 4'b0111; // x=14, y=1
        pixel_data[1][15] = 4'b0111; // x=15, y=1
        pixel_data[1][16] = 4'b0111; // x=16, y=1
        pixel_data[1][17] = 4'b0111; // x=17, y=1
        pixel_data[1][18] = 4'b0111; // x=18, y=1
        pixel_data[1][19] = 4'b0111; // x=19, y=1
        pixel_data[1][20] = 4'b0111; // x=20, y=1
        pixel_data[1][21] = 4'b0111; // x=21, y=1
        pixel_data[1][22] = 4'b0111; // x=22, y=1
        pixel_data[1][23] = 4'b0111; // x=23, y=1
        pixel_data[1][24] = 4'b0111; // x=24, y=1
        pixel_data[1][25] = 4'b0111; // x=25, y=1
        pixel_data[1][26] = 4'b0111; // x=26, y=1
        pixel_data[1][27] = 4'b0111; // x=27, y=1
        pixel_data[1][28] = 4'b0111; // x=28, y=1
        pixel_data[1][29] = 4'b0111; // x=29, y=1
        pixel_data[1][30] = 4'b0111; // x=30, y=1
        pixel_data[1][31] = 4'b0111; // x=31, y=1
        pixel_data[1][32] = 4'b0111; // x=32, y=1
        pixel_data[1][33] = 4'b0111; // x=33, y=1
        pixel_data[1][34] = 4'b0111; // x=34, y=1
        pixel_data[1][35] = 4'b0111; // x=35, y=1
        pixel_data[1][36] = 4'b0111; // x=36, y=1
        pixel_data[1][37] = 4'b0111; // x=37, y=1
        pixel_data[1][38] = 4'b0111; // x=38, y=1
        pixel_data[1][39] = 4'b0111; // x=39, y=1
        pixel_data[1][40] = 4'b0111; // x=40, y=1
        pixel_data[1][41] = 4'b0111; // x=41, y=1
        pixel_data[1][42] = 4'b0111; // x=42, y=1
        pixel_data[1][43] = 4'b0111; // x=43, y=1
        pixel_data[1][44] = 4'b0111; // x=44, y=1
        pixel_data[1][45] = 4'b0111; // x=45, y=1
        pixel_data[1][46] = 4'b0111; // x=46, y=1
        pixel_data[1][47] = 4'b0111; // x=47, y=1
        pixel_data[1][48] = 4'b0111; // x=48, y=1
        pixel_data[1][49] = 4'b0111; // x=49, y=1
        pixel_data[1][50] = 4'b0111; // x=50, y=1
        pixel_data[1][51] = 4'b0111; // x=51, y=1
        pixel_data[1][52] = 4'b0111; // x=52, y=1
        pixel_data[1][53] = 4'b0111; // x=53, y=1
        pixel_data[1][54] = 4'b0111; // x=54, y=1
        pixel_data[1][55] = 4'b0111; // x=55, y=1
        pixel_data[1][56] = 4'b0111; // x=56, y=1
        pixel_data[1][57] = 4'b0111; // x=57, y=1
        pixel_data[1][58] = 4'b0111; // x=58, y=1
        pixel_data[1][59] = 4'b0111; // x=59, y=1
        pixel_data[1][60] = 4'b0111; // x=60, y=1
        pixel_data[1][61] = 4'b0111; // x=61, y=1
        pixel_data[1][62] = 4'b0111; // x=62, y=1
        pixel_data[1][63] = 4'b0111; // x=63, y=1
        pixel_data[1][64] = 4'b0111; // x=64, y=1
        pixel_data[1][65] = 4'b0111; // x=65, y=1
        pixel_data[1][66] = 4'b0111; // x=66, y=1
        pixel_data[1][67] = 4'b0111; // x=67, y=1
        pixel_data[1][68] = 4'b0111; // x=68, y=1
        pixel_data[1][69] = 4'b0111; // x=69, y=1
        pixel_data[1][70] = 4'b0111; // x=70, y=1
        pixel_data[1][71] = 4'b0111; // x=71, y=1
        pixel_data[1][72] = 4'b0111; // x=72, y=1
        pixel_data[1][73] = 4'b0111; // x=73, y=1
        pixel_data[1][74] = 4'b0111; // x=74, y=1
        pixel_data[1][75] = 4'b0111; // x=75, y=1
        pixel_data[1][76] = 4'b0111; // x=76, y=1
        pixel_data[1][77] = 4'b0111; // x=77, y=1
        pixel_data[1][78] = 4'b0111; // x=78, y=1
        pixel_data[1][79] = 4'b0111; // x=79, y=1
        pixel_data[1][80] = 4'b0111; // x=80, y=1
        pixel_data[1][81] = 4'b0111; // x=81, y=1
        pixel_data[1][82] = 4'b0111; // x=82, y=1
        pixel_data[1][83] = 4'b0111; // x=83, y=1
        pixel_data[1][84] = 4'b0111; // x=84, y=1
        pixel_data[1][85] = 4'b0111; // x=85, y=1
        pixel_data[1][86] = 4'b0111; // x=86, y=1
        pixel_data[1][87] = 4'b0111; // x=87, y=1
        pixel_data[1][88] = 4'b0111; // x=88, y=1
        pixel_data[1][89] = 4'b0111; // x=89, y=1
        pixel_data[1][90] = 4'b0111; // x=90, y=1
        pixel_data[1][91] = 4'b0111; // x=91, y=1
        pixel_data[1][92] = 4'b0111; // x=92, y=1
        pixel_data[1][93] = 4'b0111; // x=93, y=1
        pixel_data[1][94] = 4'b0111; // x=94, y=1
        pixel_data[1][95] = 4'b0111; // x=95, y=1
        pixel_data[1][96] = 4'b0111; // x=96, y=1
        pixel_data[1][97] = 4'b0111; // x=97, y=1
        pixel_data[1][98] = 4'b0111; // x=98, y=1
        pixel_data[1][99] = 4'b0111; // x=99, y=1
        pixel_data[1][100] = 4'b0111; // x=100, y=1
        pixel_data[1][101] = 4'b0111; // x=101, y=1
        pixel_data[1][102] = 4'b0111; // x=102, y=1
        pixel_data[1][103] = 4'b0111; // x=103, y=1
        pixel_data[1][104] = 4'b0111; // x=104, y=1
        pixel_data[1][105] = 4'b0111; // x=105, y=1
        pixel_data[1][106] = 4'b0111; // x=106, y=1
        pixel_data[1][107] = 4'b0111; // x=107, y=1
        pixel_data[1][108] = 4'b0111; // x=108, y=1
        pixel_data[1][109] = 4'b0111; // x=109, y=1
        pixel_data[1][110] = 4'b0111; // x=110, y=1
        pixel_data[1][111] = 4'b0111; // x=111, y=1
        pixel_data[1][112] = 4'b0111; // x=112, y=1
        pixel_data[1][113] = 4'b0111; // x=113, y=1
        pixel_data[1][114] = 4'b0111; // x=114, y=1
        pixel_data[1][115] = 4'b0111; // x=115, y=1
        pixel_data[1][116] = 4'b0111; // x=116, y=1
        pixel_data[1][117] = 4'b0111; // x=117, y=1
        pixel_data[1][118] = 4'b0111; // x=118, y=1
        pixel_data[1][119] = 4'b0111; // x=119, y=1
        pixel_data[1][120] = 4'b0111; // x=120, y=1
        pixel_data[1][121] = 4'b0111; // x=121, y=1
        pixel_data[1][122] = 4'b0111; // x=122, y=1
        pixel_data[1][123] = 4'b0111; // x=123, y=1
        pixel_data[1][124] = 4'b0111; // x=124, y=1
        pixel_data[1][125] = 4'b0111; // x=125, y=1
        pixel_data[1][126] = 4'b0111; // x=126, y=1
        pixel_data[1][127] = 4'b0111; // x=127, y=1
        pixel_data[1][128] = 4'b0111; // x=128, y=1
        pixel_data[1][129] = 4'b0111; // x=129, y=1
        pixel_data[1][130] = 4'b0111; // x=130, y=1
        pixel_data[1][131] = 4'b0111; // x=131, y=1
        pixel_data[1][132] = 4'b0111; // x=132, y=1
        pixel_data[1][133] = 4'b0111; // x=133, y=1
        pixel_data[1][134] = 4'b0111; // x=134, y=1
        pixel_data[1][135] = 4'b0111; // x=135, y=1
        pixel_data[1][136] = 4'b0111; // x=136, y=1
        pixel_data[1][137] = 4'b0111; // x=137, y=1
        pixel_data[1][138] = 4'b0111; // x=138, y=1
        pixel_data[1][139] = 4'b0111; // x=139, y=1
        pixel_data[1][140] = 4'b0111; // x=140, y=1
        pixel_data[1][141] = 4'b0111; // x=141, y=1
        pixel_data[1][142] = 4'b0111; // x=142, y=1
        pixel_data[1][143] = 4'b0111; // x=143, y=1
        pixel_data[1][144] = 4'b0111; // x=144, y=1
        pixel_data[1][145] = 4'b0111; // x=145, y=1
        pixel_data[1][146] = 4'b0111; // x=146, y=1
        pixel_data[1][147] = 4'b0111; // x=147, y=1
        pixel_data[1][148] = 4'b0111; // x=148, y=1
        pixel_data[1][149] = 4'b0111; // x=149, y=1
        pixel_data[1][150] = 4'b0111; // x=150, y=1
        pixel_data[1][151] = 4'b0111; // x=151, y=1
        pixel_data[1][152] = 4'b0111; // x=152, y=1
        pixel_data[1][153] = 4'b0111; // x=153, y=1
        pixel_data[1][154] = 4'b0111; // x=154, y=1
        pixel_data[1][155] = 4'b0111; // x=155, y=1
        pixel_data[1][156] = 4'b0111; // x=156, y=1
        pixel_data[1][157] = 4'b0111; // x=157, y=1
        pixel_data[1][158] = 4'b0111; // x=158, y=1
        pixel_data[1][159] = 4'b0111; // x=159, y=1
        pixel_data[1][160] = 4'b0111; // x=160, y=1
        pixel_data[1][161] = 4'b0111; // x=161, y=1
        pixel_data[1][162] = 4'b0111; // x=162, y=1
        pixel_data[1][163] = 4'b0111; // x=163, y=1
        pixel_data[1][164] = 4'b0111; // x=164, y=1
        pixel_data[1][165] = 4'b0111; // x=165, y=1
        pixel_data[1][166] = 4'b0111; // x=166, y=1
        pixel_data[1][167] = 4'b0111; // x=167, y=1
        pixel_data[1][168] = 4'b0111; // x=168, y=1
        pixel_data[1][169] = 4'b0111; // x=169, y=1
        pixel_data[1][170] = 4'b0111; // x=170, y=1
        pixel_data[1][171] = 4'b0111; // x=171, y=1
        pixel_data[1][172] = 4'b0111; // x=172, y=1
        pixel_data[1][173] = 4'b0111; // x=173, y=1
        pixel_data[1][174] = 4'b0111; // x=174, y=1
        pixel_data[1][175] = 4'b0111; // x=175, y=1
        pixel_data[1][176] = 4'b0111; // x=176, y=1
        pixel_data[1][177] = 4'b0111; // x=177, y=1
        pixel_data[1][178] = 4'b0111; // x=178, y=1
        pixel_data[1][179] = 4'b0111; // x=179, y=1
        pixel_data[2][0] = 4'b0111; // x=0, y=2
        pixel_data[2][1] = 4'b0111; // x=1, y=2
        pixel_data[2][2] = 4'b0111; // x=2, y=2
        pixel_data[2][3] = 4'b0111; // x=3, y=2
        pixel_data[2][4] = 4'b0111; // x=4, y=2
        pixel_data[2][5] = 4'b0111; // x=5, y=2
        pixel_data[2][6] = 4'b0111; // x=6, y=2
        pixel_data[2][7] = 4'b0111; // x=7, y=2
        pixel_data[2][8] = 4'b0111; // x=8, y=2
        pixel_data[2][9] = 4'b0111; // x=9, y=2
        pixel_data[2][10] = 4'b0111; // x=10, y=2
        pixel_data[2][11] = 4'b0111; // x=11, y=2
        pixel_data[2][12] = 4'b0111; // x=12, y=2
        pixel_data[2][13] = 4'b0111; // x=13, y=2
        pixel_data[2][14] = 4'b0111; // x=14, y=2
        pixel_data[2][15] = 4'b0111; // x=15, y=2
        pixel_data[2][16] = 4'b0111; // x=16, y=2
        pixel_data[2][17] = 4'b0111; // x=17, y=2
        pixel_data[2][18] = 4'b0111; // x=18, y=2
        pixel_data[2][19] = 4'b0111; // x=19, y=2
        pixel_data[2][20] = 4'b0111; // x=20, y=2
        pixel_data[2][21] = 4'b0111; // x=21, y=2
        pixel_data[2][22] = 4'b0111; // x=22, y=2
        pixel_data[2][23] = 4'b0111; // x=23, y=2
        pixel_data[2][24] = 4'b0111; // x=24, y=2
        pixel_data[2][25] = 4'b0111; // x=25, y=2
        pixel_data[2][26] = 4'b0111; // x=26, y=2
        pixel_data[2][27] = 4'b0111; // x=27, y=2
        pixel_data[2][28] = 4'b0111; // x=28, y=2
        pixel_data[2][29] = 4'b0111; // x=29, y=2
        pixel_data[2][30] = 4'b0111; // x=30, y=2
        pixel_data[2][31] = 4'b0111; // x=31, y=2
        pixel_data[2][32] = 4'b0111; // x=32, y=2
        pixel_data[2][33] = 4'b0111; // x=33, y=2
        pixel_data[2][34] = 4'b0111; // x=34, y=2
        pixel_data[2][35] = 4'b0111; // x=35, y=2
        pixel_data[2][36] = 4'b0111; // x=36, y=2
        pixel_data[2][37] = 4'b0111; // x=37, y=2
        pixel_data[2][38] = 4'b0111; // x=38, y=2
        pixel_data[2][39] = 4'b0111; // x=39, y=2
        pixel_data[2][40] = 4'b0111; // x=40, y=2
        pixel_data[2][41] = 4'b0111; // x=41, y=2
        pixel_data[2][42] = 4'b0111; // x=42, y=2
        pixel_data[2][43] = 4'b0111; // x=43, y=2
        pixel_data[2][44] = 4'b0111; // x=44, y=2
        pixel_data[2][45] = 4'b0111; // x=45, y=2
        pixel_data[2][46] = 4'b0111; // x=46, y=2
        pixel_data[2][47] = 4'b0111; // x=47, y=2
        pixel_data[2][48] = 4'b0111; // x=48, y=2
        pixel_data[2][49] = 4'b0111; // x=49, y=2
        pixel_data[2][50] = 4'b0111; // x=50, y=2
        pixel_data[2][51] = 4'b0111; // x=51, y=2
        pixel_data[2][52] = 4'b0111; // x=52, y=2
        pixel_data[2][53] = 4'b0111; // x=53, y=2
        pixel_data[2][54] = 4'b0111; // x=54, y=2
        pixel_data[2][55] = 4'b0111; // x=55, y=2
        pixel_data[2][56] = 4'b0111; // x=56, y=2
        pixel_data[2][57] = 4'b0111; // x=57, y=2
        pixel_data[2][58] = 4'b0111; // x=58, y=2
        pixel_data[2][59] = 4'b0111; // x=59, y=2
        pixel_data[2][60] = 4'b0111; // x=60, y=2
        pixel_data[2][61] = 4'b0111; // x=61, y=2
        pixel_data[2][62] = 4'b0111; // x=62, y=2
        pixel_data[2][63] = 4'b0111; // x=63, y=2
        pixel_data[2][64] = 4'b0111; // x=64, y=2
        pixel_data[2][65] = 4'b0111; // x=65, y=2
        pixel_data[2][66] = 4'b0111; // x=66, y=2
        pixel_data[2][67] = 4'b0111; // x=67, y=2
        pixel_data[2][68] = 4'b0111; // x=68, y=2
        pixel_data[2][69] = 4'b0111; // x=69, y=2
        pixel_data[2][70] = 4'b0111; // x=70, y=2
        pixel_data[2][71] = 4'b0111; // x=71, y=2
        pixel_data[2][72] = 4'b0111; // x=72, y=2
        pixel_data[2][73] = 4'b0111; // x=73, y=2
        pixel_data[2][74] = 4'b0111; // x=74, y=2
        pixel_data[2][75] = 4'b0111; // x=75, y=2
        pixel_data[2][76] = 4'b0111; // x=76, y=2
        pixel_data[2][77] = 4'b0111; // x=77, y=2
        pixel_data[2][78] = 4'b0111; // x=78, y=2
        pixel_data[2][79] = 4'b0111; // x=79, y=2
        pixel_data[2][80] = 4'b0111; // x=80, y=2
        pixel_data[2][81] = 4'b0111; // x=81, y=2
        pixel_data[2][82] = 4'b0111; // x=82, y=2
        pixel_data[2][83] = 4'b0111; // x=83, y=2
        pixel_data[2][84] = 4'b0111; // x=84, y=2
        pixel_data[2][85] = 4'b0111; // x=85, y=2
        pixel_data[2][86] = 4'b0111; // x=86, y=2
        pixel_data[2][87] = 4'b0111; // x=87, y=2
        pixel_data[2][88] = 4'b0111; // x=88, y=2
        pixel_data[2][89] = 4'b0111; // x=89, y=2
        pixel_data[2][90] = 4'b0111; // x=90, y=2
        pixel_data[2][91] = 4'b0111; // x=91, y=2
        pixel_data[2][92] = 4'b0111; // x=92, y=2
        pixel_data[2][93] = 4'b0111; // x=93, y=2
        pixel_data[2][94] = 4'b0111; // x=94, y=2
        pixel_data[2][95] = 4'b0111; // x=95, y=2
        pixel_data[2][96] = 4'b0111; // x=96, y=2
        pixel_data[2][97] = 4'b0111; // x=97, y=2
        pixel_data[2][98] = 4'b0111; // x=98, y=2
        pixel_data[2][99] = 4'b0111; // x=99, y=2
        pixel_data[2][100] = 4'b0111; // x=100, y=2
        pixel_data[2][101] = 4'b0111; // x=101, y=2
        pixel_data[2][102] = 4'b0111; // x=102, y=2
        pixel_data[2][103] = 4'b0111; // x=103, y=2
        pixel_data[2][104] = 4'b0111; // x=104, y=2
        pixel_data[2][105] = 4'b0111; // x=105, y=2
        pixel_data[2][106] = 4'b0111; // x=106, y=2
        pixel_data[2][107] = 4'b0111; // x=107, y=2
        pixel_data[2][108] = 4'b0111; // x=108, y=2
        pixel_data[2][109] = 4'b0111; // x=109, y=2
        pixel_data[2][110] = 4'b0111; // x=110, y=2
        pixel_data[2][111] = 4'b0111; // x=111, y=2
        pixel_data[2][112] = 4'b0111; // x=112, y=2
        pixel_data[2][113] = 4'b0111; // x=113, y=2
        pixel_data[2][114] = 4'b0111; // x=114, y=2
        pixel_data[2][115] = 4'b0111; // x=115, y=2
        pixel_data[2][116] = 4'b0111; // x=116, y=2
        pixel_data[2][117] = 4'b0111; // x=117, y=2
        pixel_data[2][118] = 4'b0111; // x=118, y=2
        pixel_data[2][119] = 4'b0111; // x=119, y=2
        pixel_data[2][120] = 4'b0111; // x=120, y=2
        pixel_data[2][121] = 4'b0111; // x=121, y=2
        pixel_data[2][122] = 4'b0111; // x=122, y=2
        pixel_data[2][123] = 4'b0111; // x=123, y=2
        pixel_data[2][124] = 4'b0111; // x=124, y=2
        pixel_data[2][125] = 4'b0111; // x=125, y=2
        pixel_data[2][126] = 4'b0111; // x=126, y=2
        pixel_data[2][127] = 4'b0111; // x=127, y=2
        pixel_data[2][128] = 4'b0111; // x=128, y=2
        pixel_data[2][129] = 4'b0111; // x=129, y=2
        pixel_data[2][130] = 4'b0111; // x=130, y=2
        pixel_data[2][131] = 4'b0111; // x=131, y=2
        pixel_data[2][132] = 4'b0111; // x=132, y=2
        pixel_data[2][133] = 4'b0111; // x=133, y=2
        pixel_data[2][134] = 4'b0111; // x=134, y=2
        pixel_data[2][135] = 4'b0111; // x=135, y=2
        pixel_data[2][136] = 4'b0111; // x=136, y=2
        pixel_data[2][137] = 4'b0111; // x=137, y=2
        pixel_data[2][138] = 4'b0111; // x=138, y=2
        pixel_data[2][139] = 4'b0111; // x=139, y=2
        pixel_data[2][140] = 4'b0111; // x=140, y=2
        pixel_data[2][141] = 4'b0111; // x=141, y=2
        pixel_data[2][142] = 4'b0111; // x=142, y=2
        pixel_data[2][143] = 4'b0111; // x=143, y=2
        pixel_data[2][144] = 4'b0111; // x=144, y=2
        pixel_data[2][145] = 4'b0111; // x=145, y=2
        pixel_data[2][146] = 4'b0111; // x=146, y=2
        pixel_data[2][147] = 4'b0111; // x=147, y=2
        pixel_data[2][148] = 4'b0111; // x=148, y=2
        pixel_data[2][149] = 4'b0111; // x=149, y=2
        pixel_data[2][150] = 4'b0111; // x=150, y=2
        pixel_data[2][151] = 4'b0111; // x=151, y=2
        pixel_data[2][152] = 4'b0111; // x=152, y=2
        pixel_data[2][153] = 4'b0111; // x=153, y=2
        pixel_data[2][154] = 4'b0111; // x=154, y=2
        pixel_data[2][155] = 4'b0111; // x=155, y=2
        pixel_data[2][156] = 4'b0111; // x=156, y=2
        pixel_data[2][157] = 4'b0111; // x=157, y=2
        pixel_data[2][158] = 4'b0111; // x=158, y=2
        pixel_data[2][159] = 4'b0111; // x=159, y=2
        pixel_data[2][160] = 4'b0111; // x=160, y=2
        pixel_data[2][161] = 4'b0111; // x=161, y=2
        pixel_data[2][162] = 4'b0111; // x=162, y=2
        pixel_data[2][163] = 4'b0111; // x=163, y=2
        pixel_data[2][164] = 4'b0111; // x=164, y=2
        pixel_data[2][165] = 4'b0111; // x=165, y=2
        pixel_data[2][166] = 4'b0111; // x=166, y=2
        pixel_data[2][167] = 4'b0111; // x=167, y=2
        pixel_data[2][168] = 4'b0111; // x=168, y=2
        pixel_data[2][169] = 4'b0111; // x=169, y=2
        pixel_data[2][170] = 4'b0111; // x=170, y=2
        pixel_data[2][171] = 4'b0111; // x=171, y=2
        pixel_data[2][172] = 4'b0111; // x=172, y=2
        pixel_data[2][173] = 4'b0111; // x=173, y=2
        pixel_data[2][174] = 4'b0111; // x=174, y=2
        pixel_data[2][175] = 4'b0111; // x=175, y=2
        pixel_data[2][176] = 4'b0111; // x=176, y=2
        pixel_data[2][177] = 4'b0111; // x=177, y=2
        pixel_data[2][178] = 4'b0111; // x=178, y=2
        pixel_data[2][179] = 4'b0111; // x=179, y=2
        pixel_data[3][0] = 4'b0111; // x=0, y=3
        pixel_data[3][1] = 4'b0111; // x=1, y=3
        pixel_data[3][2] = 4'b0111; // x=2, y=3
        pixel_data[3][3] = 4'b0111; // x=3, y=3
        pixel_data[3][4] = 4'b0111; // x=4, y=3
        pixel_data[3][5] = 4'b0111; // x=5, y=3
        pixel_data[3][6] = 4'b0111; // x=6, y=3
        pixel_data[3][7] = 4'b0111; // x=7, y=3
        pixel_data[3][8] = 4'b0111; // x=8, y=3
        pixel_data[3][9] = 4'b0111; // x=9, y=3
        pixel_data[3][10] = 4'b0111; // x=10, y=3
        pixel_data[3][11] = 4'b0111; // x=11, y=3
        pixel_data[3][12] = 4'b0111; // x=12, y=3
        pixel_data[3][13] = 4'b0111; // x=13, y=3
        pixel_data[3][14] = 4'b0111; // x=14, y=3
        pixel_data[3][15] = 4'b0111; // x=15, y=3
        pixel_data[3][16] = 4'b0111; // x=16, y=3
        pixel_data[3][17] = 4'b0111; // x=17, y=3
        pixel_data[3][18] = 4'b0111; // x=18, y=3
        pixel_data[3][19] = 4'b0111; // x=19, y=3
        pixel_data[3][20] = 4'b0111; // x=20, y=3
        pixel_data[3][21] = 4'b0111; // x=21, y=3
        pixel_data[3][22] = 4'b0111; // x=22, y=3
        pixel_data[3][23] = 4'b0111; // x=23, y=3
        pixel_data[3][24] = 4'b0111; // x=24, y=3
        pixel_data[3][25] = 4'b0111; // x=25, y=3
        pixel_data[3][26] = 4'b0111; // x=26, y=3
        pixel_data[3][27] = 4'b0111; // x=27, y=3
        pixel_data[3][28] = 4'b0111; // x=28, y=3
        pixel_data[3][29] = 4'b0111; // x=29, y=3
        pixel_data[3][30] = 4'b0111; // x=30, y=3
        pixel_data[3][31] = 4'b0111; // x=31, y=3
        pixel_data[3][32] = 4'b0111; // x=32, y=3
        pixel_data[3][33] = 4'b0111; // x=33, y=3
        pixel_data[3][34] = 4'b0111; // x=34, y=3
        pixel_data[3][35] = 4'b0111; // x=35, y=3
        pixel_data[3][36] = 4'b0111; // x=36, y=3
        pixel_data[3][37] = 4'b0111; // x=37, y=3
        pixel_data[3][38] = 4'b0111; // x=38, y=3
        pixel_data[3][39] = 4'b0111; // x=39, y=3
        pixel_data[3][40] = 4'b0111; // x=40, y=3
        pixel_data[3][41] = 4'b0111; // x=41, y=3
        pixel_data[3][42] = 4'b0111; // x=42, y=3
        pixel_data[3][43] = 4'b0111; // x=43, y=3
        pixel_data[3][44] = 4'b0111; // x=44, y=3
        pixel_data[3][45] = 4'b0111; // x=45, y=3
        pixel_data[3][46] = 4'b0111; // x=46, y=3
        pixel_data[3][47] = 4'b0111; // x=47, y=3
        pixel_data[3][48] = 4'b0111; // x=48, y=3
        pixel_data[3][49] = 4'b0111; // x=49, y=3
        pixel_data[3][50] = 4'b0111; // x=50, y=3
        pixel_data[3][51] = 4'b0111; // x=51, y=3
        pixel_data[3][52] = 4'b0111; // x=52, y=3
        pixel_data[3][53] = 4'b0111; // x=53, y=3
        pixel_data[3][54] = 4'b0111; // x=54, y=3
        pixel_data[3][55] = 4'b0111; // x=55, y=3
        pixel_data[3][56] = 4'b0111; // x=56, y=3
        pixel_data[3][57] = 4'b0111; // x=57, y=3
        pixel_data[3][58] = 4'b0111; // x=58, y=3
        pixel_data[3][59] = 4'b0111; // x=59, y=3
        pixel_data[3][60] = 4'b0111; // x=60, y=3
        pixel_data[3][61] = 4'b0111; // x=61, y=3
        pixel_data[3][62] = 4'b0111; // x=62, y=3
        pixel_data[3][63] = 4'b0111; // x=63, y=3
        pixel_data[3][64] = 4'b0111; // x=64, y=3
        pixel_data[3][65] = 4'b0111; // x=65, y=3
        pixel_data[3][66] = 4'b0111; // x=66, y=3
        pixel_data[3][67] = 4'b0111; // x=67, y=3
        pixel_data[3][68] = 4'b0111; // x=68, y=3
        pixel_data[3][69] = 4'b0111; // x=69, y=3
        pixel_data[3][70] = 4'b0111; // x=70, y=3
        pixel_data[3][71] = 4'b0111; // x=71, y=3
        pixel_data[3][72] = 4'b0111; // x=72, y=3
        pixel_data[3][73] = 4'b0111; // x=73, y=3
        pixel_data[3][74] = 4'b0111; // x=74, y=3
        pixel_data[3][75] = 4'b0111; // x=75, y=3
        pixel_data[3][76] = 4'b0111; // x=76, y=3
        pixel_data[3][77] = 4'b0111; // x=77, y=3
        pixel_data[3][78] = 4'b0111; // x=78, y=3
        pixel_data[3][79] = 4'b0111; // x=79, y=3
        pixel_data[3][80] = 4'b0111; // x=80, y=3
        pixel_data[3][81] = 4'b0111; // x=81, y=3
        pixel_data[3][82] = 4'b0111; // x=82, y=3
        pixel_data[3][83] = 4'b0111; // x=83, y=3
        pixel_data[3][84] = 4'b0111; // x=84, y=3
        pixel_data[3][85] = 4'b0111; // x=85, y=3
        pixel_data[3][86] = 4'b0111; // x=86, y=3
        pixel_data[3][87] = 4'b0111; // x=87, y=3
        pixel_data[3][88] = 4'b0111; // x=88, y=3
        pixel_data[3][89] = 4'b0111; // x=89, y=3
        pixel_data[3][90] = 4'b0111; // x=90, y=3
        pixel_data[3][91] = 4'b0111; // x=91, y=3
        pixel_data[3][92] = 4'b0111; // x=92, y=3
        pixel_data[3][93] = 4'b0111; // x=93, y=3
        pixel_data[3][94] = 4'b0111; // x=94, y=3
        pixel_data[3][95] = 4'b0111; // x=95, y=3
        pixel_data[3][96] = 4'b0111; // x=96, y=3
        pixel_data[3][97] = 4'b0111; // x=97, y=3
        pixel_data[3][98] = 4'b0111; // x=98, y=3
        pixel_data[3][99] = 4'b0111; // x=99, y=3
        pixel_data[3][100] = 4'b0111; // x=100, y=3
        pixel_data[3][101] = 4'b0111; // x=101, y=3
        pixel_data[3][102] = 4'b0111; // x=102, y=3
        pixel_data[3][103] = 4'b0111; // x=103, y=3
        pixel_data[3][104] = 4'b0111; // x=104, y=3
        pixel_data[3][105] = 4'b0111; // x=105, y=3
        pixel_data[3][106] = 4'b0111; // x=106, y=3
        pixel_data[3][107] = 4'b0111; // x=107, y=3
        pixel_data[3][108] = 4'b0111; // x=108, y=3
        pixel_data[3][109] = 4'b0111; // x=109, y=3
        pixel_data[3][110] = 4'b0111; // x=110, y=3
        pixel_data[3][111] = 4'b0111; // x=111, y=3
        pixel_data[3][112] = 4'b0111; // x=112, y=3
        pixel_data[3][113] = 4'b0111; // x=113, y=3
        pixel_data[3][114] = 4'b0111; // x=114, y=3
        pixel_data[3][115] = 4'b0111; // x=115, y=3
        pixel_data[3][116] = 4'b0111; // x=116, y=3
        pixel_data[3][117] = 4'b0111; // x=117, y=3
        pixel_data[3][118] = 4'b0111; // x=118, y=3
        pixel_data[3][119] = 4'b0111; // x=119, y=3
        pixel_data[3][120] = 4'b0111; // x=120, y=3
        pixel_data[3][121] = 4'b0111; // x=121, y=3
        pixel_data[3][122] = 4'b0111; // x=122, y=3
        pixel_data[3][123] = 4'b0111; // x=123, y=3
        pixel_data[3][124] = 4'b0111; // x=124, y=3
        pixel_data[3][125] = 4'b0111; // x=125, y=3
        pixel_data[3][126] = 4'b0111; // x=126, y=3
        pixel_data[3][127] = 4'b0111; // x=127, y=3
        pixel_data[3][128] = 4'b0111; // x=128, y=3
        pixel_data[3][129] = 4'b0111; // x=129, y=3
        pixel_data[3][130] = 4'b0111; // x=130, y=3
        pixel_data[3][131] = 4'b0111; // x=131, y=3
        pixel_data[3][132] = 4'b0111; // x=132, y=3
        pixel_data[3][133] = 4'b0111; // x=133, y=3
        pixel_data[3][134] = 4'b0111; // x=134, y=3
        pixel_data[3][135] = 4'b0111; // x=135, y=3
        pixel_data[3][136] = 4'b0111; // x=136, y=3
        pixel_data[3][137] = 4'b0111; // x=137, y=3
        pixel_data[3][138] = 4'b0111; // x=138, y=3
        pixel_data[3][139] = 4'b0111; // x=139, y=3
        pixel_data[3][140] = 4'b0111; // x=140, y=3
        pixel_data[3][141] = 4'b0111; // x=141, y=3
        pixel_data[3][142] = 4'b0111; // x=142, y=3
        pixel_data[3][143] = 4'b0111; // x=143, y=3
        pixel_data[3][144] = 4'b0111; // x=144, y=3
        pixel_data[3][145] = 4'b0111; // x=145, y=3
        pixel_data[3][146] = 4'b0111; // x=146, y=3
        pixel_data[3][147] = 4'b0111; // x=147, y=3
        pixel_data[3][148] = 4'b0111; // x=148, y=3
        pixel_data[3][149] = 4'b0111; // x=149, y=3
        pixel_data[3][150] = 4'b0111; // x=150, y=3
        pixel_data[3][151] = 4'b0111; // x=151, y=3
        pixel_data[3][152] = 4'b0111; // x=152, y=3
        pixel_data[3][153] = 4'b0111; // x=153, y=3
        pixel_data[3][154] = 4'b0111; // x=154, y=3
        pixel_data[3][155] = 4'b0111; // x=155, y=3
        pixel_data[3][156] = 4'b0111; // x=156, y=3
        pixel_data[3][157] = 4'b0111; // x=157, y=3
        pixel_data[3][158] = 4'b0111; // x=158, y=3
        pixel_data[3][159] = 4'b0111; // x=159, y=3
        pixel_data[3][160] = 4'b0111; // x=160, y=3
        pixel_data[3][161] = 4'b0111; // x=161, y=3
        pixel_data[3][162] = 4'b0111; // x=162, y=3
        pixel_data[3][163] = 4'b0111; // x=163, y=3
        pixel_data[3][164] = 4'b0111; // x=164, y=3
        pixel_data[3][165] = 4'b0111; // x=165, y=3
        pixel_data[3][166] = 4'b0111; // x=166, y=3
        pixel_data[3][167] = 4'b0111; // x=167, y=3
        pixel_data[3][168] = 4'b0111; // x=168, y=3
        pixel_data[3][169] = 4'b0111; // x=169, y=3
        pixel_data[3][170] = 4'b0111; // x=170, y=3
        pixel_data[3][171] = 4'b0111; // x=171, y=3
        pixel_data[3][172] = 4'b0111; // x=172, y=3
        pixel_data[3][173] = 4'b0111; // x=173, y=3
        pixel_data[3][174] = 4'b0111; // x=174, y=3
        pixel_data[3][175] = 4'b0111; // x=175, y=3
        pixel_data[3][176] = 4'b0111; // x=176, y=3
        pixel_data[3][177] = 4'b0111; // x=177, y=3
        pixel_data[3][178] = 4'b0111; // x=178, y=3
        pixel_data[3][179] = 4'b0111; // x=179, y=3
        pixel_data[4][0] = 4'b0111; // x=0, y=4
        pixel_data[4][1] = 4'b0111; // x=1, y=4
        pixel_data[4][2] = 4'b0111; // x=2, y=4
        pixel_data[4][3] = 4'b0111; // x=3, y=4
        pixel_data[4][4] = 4'b0111; // x=4, y=4
        pixel_data[4][5] = 4'b0111; // x=5, y=4
        pixel_data[4][6] = 4'b0111; // x=6, y=4
        pixel_data[4][7] = 4'b0111; // x=7, y=4
        pixel_data[4][8] = 4'b0111; // x=8, y=4
        pixel_data[4][9] = 4'b0111; // x=9, y=4
        pixel_data[4][10] = 4'b0111; // x=10, y=4
        pixel_data[4][11] = 4'b0111; // x=11, y=4
        pixel_data[4][12] = 4'b0111; // x=12, y=4
        pixel_data[4][13] = 4'b0111; // x=13, y=4
        pixel_data[4][14] = 4'b0111; // x=14, y=4
        pixel_data[4][15] = 4'b0111; // x=15, y=4
        pixel_data[4][16] = 4'b0111; // x=16, y=4
        pixel_data[4][17] = 4'b0111; // x=17, y=4
        pixel_data[4][18] = 4'b0111; // x=18, y=4
        pixel_data[4][19] = 4'b0111; // x=19, y=4
        pixel_data[4][20] = 4'b0111; // x=20, y=4
        pixel_data[4][21] = 4'b0111; // x=21, y=4
        pixel_data[4][22] = 4'b0111; // x=22, y=4
        pixel_data[4][23] = 4'b0111; // x=23, y=4
        pixel_data[4][24] = 4'b0111; // x=24, y=4
        pixel_data[4][25] = 4'b0111; // x=25, y=4
        pixel_data[4][26] = 4'b0111; // x=26, y=4
        pixel_data[4][27] = 4'b0111; // x=27, y=4
        pixel_data[4][28] = 4'b0111; // x=28, y=4
        pixel_data[4][29] = 4'b0111; // x=29, y=4
        pixel_data[4][30] = 4'b0111; // x=30, y=4
        pixel_data[4][31] = 4'b0111; // x=31, y=4
        pixel_data[4][32] = 4'b0111; // x=32, y=4
        pixel_data[4][33] = 4'b0111; // x=33, y=4
        pixel_data[4][34] = 4'b0111; // x=34, y=4
        pixel_data[4][35] = 4'b0111; // x=35, y=4
        pixel_data[4][36] = 4'b0111; // x=36, y=4
        pixel_data[4][37] = 4'b0111; // x=37, y=4
        pixel_data[4][38] = 4'b0111; // x=38, y=4
        pixel_data[4][39] = 4'b0111; // x=39, y=4
        pixel_data[4][40] = 4'b0111; // x=40, y=4
        pixel_data[4][41] = 4'b0111; // x=41, y=4
        pixel_data[4][42] = 4'b0111; // x=42, y=4
        pixel_data[4][43] = 4'b0111; // x=43, y=4
        pixel_data[4][44] = 4'b0111; // x=44, y=4
        pixel_data[4][45] = 4'b0111; // x=45, y=4
        pixel_data[4][46] = 4'b0111; // x=46, y=4
        pixel_data[4][47] = 4'b0111; // x=47, y=4
        pixel_data[4][48] = 4'b0111; // x=48, y=4
        pixel_data[4][49] = 4'b0111; // x=49, y=4
        pixel_data[4][50] = 4'b0111; // x=50, y=4
        pixel_data[4][51] = 4'b0111; // x=51, y=4
        pixel_data[4][52] = 4'b0111; // x=52, y=4
        pixel_data[4][53] = 4'b0111; // x=53, y=4
        pixel_data[4][54] = 4'b0111; // x=54, y=4
        pixel_data[4][55] = 4'b0111; // x=55, y=4
        pixel_data[4][56] = 4'b0111; // x=56, y=4
        pixel_data[4][57] = 4'b0111; // x=57, y=4
        pixel_data[4][58] = 4'b0111; // x=58, y=4
        pixel_data[4][59] = 4'b0111; // x=59, y=4
        pixel_data[4][60] = 4'b0111; // x=60, y=4
        pixel_data[4][61] = 4'b0111; // x=61, y=4
        pixel_data[4][62] = 4'b0111; // x=62, y=4
        pixel_data[4][63] = 4'b0111; // x=63, y=4
        pixel_data[4][64] = 4'b0111; // x=64, y=4
        pixel_data[4][65] = 4'b0111; // x=65, y=4
        pixel_data[4][66] = 4'b0111; // x=66, y=4
        pixel_data[4][67] = 4'b0111; // x=67, y=4
        pixel_data[4][68] = 4'b0111; // x=68, y=4
        pixel_data[4][69] = 4'b0111; // x=69, y=4
        pixel_data[4][70] = 4'b0111; // x=70, y=4
        pixel_data[4][71] = 4'b0111; // x=71, y=4
        pixel_data[4][72] = 4'b0111; // x=72, y=4
        pixel_data[4][73] = 4'b0111; // x=73, y=4
        pixel_data[4][74] = 4'b0111; // x=74, y=4
        pixel_data[4][75] = 4'b0111; // x=75, y=4
        pixel_data[4][76] = 4'b0111; // x=76, y=4
        pixel_data[4][77] = 4'b0111; // x=77, y=4
        pixel_data[4][78] = 4'b0111; // x=78, y=4
        pixel_data[4][79] = 4'b0111; // x=79, y=4
        pixel_data[4][80] = 4'b0111; // x=80, y=4
        pixel_data[4][81] = 4'b0111; // x=81, y=4
        pixel_data[4][82] = 4'b0111; // x=82, y=4
        pixel_data[4][83] = 4'b0111; // x=83, y=4
        pixel_data[4][84] = 4'b0111; // x=84, y=4
        pixel_data[4][85] = 4'b0111; // x=85, y=4
        pixel_data[4][86] = 4'b0111; // x=86, y=4
        pixel_data[4][87] = 4'b0111; // x=87, y=4
        pixel_data[4][88] = 4'b0111; // x=88, y=4
        pixel_data[4][89] = 4'b0111; // x=89, y=4
        pixel_data[4][90] = 4'b0111; // x=90, y=4
        pixel_data[4][91] = 4'b0111; // x=91, y=4
        pixel_data[4][92] = 4'b0111; // x=92, y=4
        pixel_data[4][93] = 4'b0111; // x=93, y=4
        pixel_data[4][94] = 4'b0111; // x=94, y=4
        pixel_data[4][95] = 4'b0111; // x=95, y=4
        pixel_data[4][96] = 4'b0111; // x=96, y=4
        pixel_data[4][97] = 4'b0111; // x=97, y=4
        pixel_data[4][98] = 4'b0111; // x=98, y=4
        pixel_data[4][99] = 4'b0111; // x=99, y=4
        pixel_data[4][100] = 4'b0111; // x=100, y=4
        pixel_data[4][101] = 4'b0111; // x=101, y=4
        pixel_data[4][102] = 4'b0111; // x=102, y=4
        pixel_data[4][103] = 4'b0111; // x=103, y=4
        pixel_data[4][104] = 4'b0111; // x=104, y=4
        pixel_data[4][105] = 4'b0111; // x=105, y=4
        pixel_data[4][106] = 4'b0111; // x=106, y=4
        pixel_data[4][107] = 4'b0111; // x=107, y=4
        pixel_data[4][108] = 4'b0111; // x=108, y=4
        pixel_data[4][109] = 4'b0111; // x=109, y=4
        pixel_data[4][110] = 4'b0111; // x=110, y=4
        pixel_data[4][111] = 4'b0111; // x=111, y=4
        pixel_data[4][112] = 4'b0111; // x=112, y=4
        pixel_data[4][113] = 4'b0111; // x=113, y=4
        pixel_data[4][114] = 4'b0111; // x=114, y=4
        pixel_data[4][115] = 4'b0111; // x=115, y=4
        pixel_data[4][116] = 4'b0111; // x=116, y=4
        pixel_data[4][117] = 4'b0111; // x=117, y=4
        pixel_data[4][118] = 4'b0111; // x=118, y=4
        pixel_data[4][119] = 4'b0111; // x=119, y=4
        pixel_data[4][120] = 4'b0111; // x=120, y=4
        pixel_data[4][121] = 4'b0111; // x=121, y=4
        pixel_data[4][122] = 4'b0111; // x=122, y=4
        pixel_data[4][123] = 4'b0111; // x=123, y=4
        pixel_data[4][124] = 4'b0111; // x=124, y=4
        pixel_data[4][125] = 4'b0111; // x=125, y=4
        pixel_data[4][126] = 4'b0111; // x=126, y=4
        pixel_data[4][127] = 4'b0111; // x=127, y=4
        pixel_data[4][128] = 4'b0111; // x=128, y=4
        pixel_data[4][129] = 4'b0111; // x=129, y=4
        pixel_data[4][130] = 4'b0111; // x=130, y=4
        pixel_data[4][131] = 4'b0111; // x=131, y=4
        pixel_data[4][132] = 4'b0111; // x=132, y=4
        pixel_data[4][133] = 4'b0111; // x=133, y=4
        pixel_data[4][134] = 4'b0111; // x=134, y=4
        pixel_data[4][135] = 4'b0111; // x=135, y=4
        pixel_data[4][136] = 4'b0111; // x=136, y=4
        pixel_data[4][137] = 4'b0111; // x=137, y=4
        pixel_data[4][138] = 4'b0111; // x=138, y=4
        pixel_data[4][139] = 4'b0111; // x=139, y=4
        pixel_data[4][140] = 4'b0111; // x=140, y=4
        pixel_data[4][141] = 4'b0111; // x=141, y=4
        pixel_data[4][142] = 4'b0111; // x=142, y=4
        pixel_data[4][143] = 4'b0111; // x=143, y=4
        pixel_data[4][144] = 4'b0111; // x=144, y=4
        pixel_data[4][145] = 4'b0111; // x=145, y=4
        pixel_data[4][146] = 4'b0111; // x=146, y=4
        pixel_data[4][147] = 4'b0111; // x=147, y=4
        pixel_data[4][148] = 4'b0111; // x=148, y=4
        pixel_data[4][149] = 4'b0111; // x=149, y=4
        pixel_data[4][150] = 4'b0111; // x=150, y=4
        pixel_data[4][151] = 4'b0111; // x=151, y=4
        pixel_data[4][152] = 4'b0111; // x=152, y=4
        pixel_data[4][153] = 4'b0111; // x=153, y=4
        pixel_data[4][154] = 4'b0111; // x=154, y=4
        pixel_data[4][155] = 4'b0111; // x=155, y=4
        pixel_data[4][156] = 4'b0111; // x=156, y=4
        pixel_data[4][157] = 4'b0111; // x=157, y=4
        pixel_data[4][158] = 4'b0111; // x=158, y=4
        pixel_data[4][159] = 4'b0111; // x=159, y=4
        pixel_data[4][160] = 4'b0111; // x=160, y=4
        pixel_data[4][161] = 4'b0111; // x=161, y=4
        pixel_data[4][162] = 4'b0111; // x=162, y=4
        pixel_data[4][163] = 4'b0111; // x=163, y=4
        pixel_data[4][164] = 4'b0111; // x=164, y=4
        pixel_data[4][165] = 4'b0111; // x=165, y=4
        pixel_data[4][166] = 4'b0111; // x=166, y=4
        pixel_data[4][167] = 4'b0111; // x=167, y=4
        pixel_data[4][168] = 4'b0111; // x=168, y=4
        pixel_data[4][169] = 4'b0111; // x=169, y=4
        pixel_data[4][170] = 4'b0111; // x=170, y=4
        pixel_data[4][171] = 4'b0111; // x=171, y=4
        pixel_data[4][172] = 4'b0111; // x=172, y=4
        pixel_data[4][173] = 4'b0111; // x=173, y=4
        pixel_data[4][174] = 4'b0111; // x=174, y=4
        pixel_data[4][175] = 4'b0111; // x=175, y=4
        pixel_data[4][176] = 4'b0111; // x=176, y=4
        pixel_data[4][177] = 4'b0111; // x=177, y=4
        pixel_data[4][178] = 4'b0111; // x=178, y=4
        pixel_data[4][179] = 4'b0111; // x=179, y=4
        pixel_data[5][0] = 4'b0111; // x=0, y=5
        pixel_data[5][1] = 4'b0111; // x=1, y=5
        pixel_data[5][2] = 4'b0111; // x=2, y=5
        pixel_data[5][3] = 4'b0111; // x=3, y=5
        pixel_data[5][4] = 4'b0111; // x=4, y=5
        pixel_data[5][5] = 4'b0111; // x=5, y=5
        pixel_data[5][6] = 4'b0111; // x=6, y=5
        pixel_data[5][7] = 4'b0111; // x=7, y=5
        pixel_data[5][8] = 4'b0111; // x=8, y=5
        pixel_data[5][9] = 4'b0111; // x=9, y=5
        pixel_data[5][10] = 4'b0111; // x=10, y=5
        pixel_data[5][11] = 4'b0111; // x=11, y=5
        pixel_data[5][12] = 4'b0111; // x=12, y=5
        pixel_data[5][13] = 4'b0111; // x=13, y=5
        pixel_data[5][14] = 4'b0111; // x=14, y=5
        pixel_data[5][15] = 4'b0111; // x=15, y=5
        pixel_data[5][16] = 4'b0111; // x=16, y=5
        pixel_data[5][17] = 4'b0111; // x=17, y=5
        pixel_data[5][18] = 4'b0111; // x=18, y=5
        pixel_data[5][19] = 4'b0111; // x=19, y=5
        pixel_data[5][20] = 4'b0111; // x=20, y=5
        pixel_data[5][21] = 4'b0111; // x=21, y=5
        pixel_data[5][22] = 4'b0111; // x=22, y=5
        pixel_data[5][23] = 4'b0111; // x=23, y=5
        pixel_data[5][24] = 4'b0111; // x=24, y=5
        pixel_data[5][25] = 4'b0111; // x=25, y=5
        pixel_data[5][26] = 4'b0111; // x=26, y=5
        pixel_data[5][27] = 4'b0111; // x=27, y=5
        pixel_data[5][28] = 4'b0111; // x=28, y=5
        pixel_data[5][29] = 4'b0111; // x=29, y=5
        pixel_data[5][30] = 4'b0111; // x=30, y=5
        pixel_data[5][31] = 4'b0111; // x=31, y=5
        pixel_data[5][32] = 4'b0111; // x=32, y=5
        pixel_data[5][33] = 4'b0111; // x=33, y=5
        pixel_data[5][34] = 4'b0111; // x=34, y=5
        pixel_data[5][35] = 4'b0111; // x=35, y=5
        pixel_data[5][36] = 4'b0111; // x=36, y=5
        pixel_data[5][37] = 4'b0111; // x=37, y=5
        pixel_data[5][38] = 4'b0111; // x=38, y=5
        pixel_data[5][39] = 4'b0111; // x=39, y=5
        pixel_data[5][40] = 4'b0111; // x=40, y=5
        pixel_data[5][41] = 4'b0111; // x=41, y=5
        pixel_data[5][42] = 4'b0111; // x=42, y=5
        pixel_data[5][43] = 4'b0111; // x=43, y=5
        pixel_data[5][44] = 4'b0111; // x=44, y=5
        pixel_data[5][45] = 4'b0111; // x=45, y=5
        pixel_data[5][46] = 4'b0111; // x=46, y=5
        pixel_data[5][47] = 4'b0111; // x=47, y=5
        pixel_data[5][48] = 4'b0111; // x=48, y=5
        pixel_data[5][49] = 4'b0111; // x=49, y=5
        pixel_data[5][50] = 4'b0111; // x=50, y=5
        pixel_data[5][51] = 4'b0111; // x=51, y=5
        pixel_data[5][52] = 4'b0111; // x=52, y=5
        pixel_data[5][53] = 4'b0111; // x=53, y=5
        pixel_data[5][54] = 4'b0111; // x=54, y=5
        pixel_data[5][55] = 4'b0111; // x=55, y=5
        pixel_data[5][56] = 4'b0111; // x=56, y=5
        pixel_data[5][57] = 4'b0111; // x=57, y=5
        pixel_data[5][58] = 4'b0111; // x=58, y=5
        pixel_data[5][59] = 4'b0111; // x=59, y=5
        pixel_data[5][60] = 4'b0111; // x=60, y=5
        pixel_data[5][61] = 4'b0111; // x=61, y=5
        pixel_data[5][62] = 4'b0111; // x=62, y=5
        pixel_data[5][63] = 4'b0111; // x=63, y=5
        pixel_data[5][64] = 4'b0111; // x=64, y=5
        pixel_data[5][65] = 4'b0111; // x=65, y=5
        pixel_data[5][66] = 4'b0111; // x=66, y=5
        pixel_data[5][67] = 4'b0111; // x=67, y=5
        pixel_data[5][68] = 4'b0111; // x=68, y=5
        pixel_data[5][69] = 4'b0111; // x=69, y=5
        pixel_data[5][70] = 4'b0111; // x=70, y=5
        pixel_data[5][71] = 4'b0111; // x=71, y=5
        pixel_data[5][72] = 4'b0111; // x=72, y=5
        pixel_data[5][73] = 4'b0111; // x=73, y=5
        pixel_data[5][74] = 4'b0111; // x=74, y=5
        pixel_data[5][75] = 4'b0111; // x=75, y=5
        pixel_data[5][76] = 4'b0111; // x=76, y=5
        pixel_data[5][77] = 4'b0111; // x=77, y=5
        pixel_data[5][78] = 4'b0111; // x=78, y=5
        pixel_data[5][79] = 4'b0111; // x=79, y=5
        pixel_data[5][80] = 4'b0111; // x=80, y=5
        pixel_data[5][81] = 4'b0111; // x=81, y=5
        pixel_data[5][82] = 4'b0111; // x=82, y=5
        pixel_data[5][83] = 4'b0111; // x=83, y=5
        pixel_data[5][84] = 4'b0111; // x=84, y=5
        pixel_data[5][85] = 4'b0111; // x=85, y=5
        pixel_data[5][86] = 4'b0111; // x=86, y=5
        pixel_data[5][87] = 4'b0111; // x=87, y=5
        pixel_data[5][88] = 4'b0111; // x=88, y=5
        pixel_data[5][89] = 4'b0111; // x=89, y=5
        pixel_data[5][90] = 4'b0111; // x=90, y=5
        pixel_data[5][91] = 4'b0111; // x=91, y=5
        pixel_data[5][92] = 4'b0111; // x=92, y=5
        pixel_data[5][93] = 4'b0111; // x=93, y=5
        pixel_data[5][94] = 4'b0111; // x=94, y=5
        pixel_data[5][95] = 4'b0111; // x=95, y=5
        pixel_data[5][96] = 4'b0111; // x=96, y=5
        pixel_data[5][97] = 4'b0111; // x=97, y=5
        pixel_data[5][98] = 4'b0111; // x=98, y=5
        pixel_data[5][99] = 4'b0111; // x=99, y=5
        pixel_data[5][100] = 4'b0111; // x=100, y=5
        pixel_data[5][101] = 4'b0111; // x=101, y=5
        pixel_data[5][102] = 4'b0111; // x=102, y=5
        pixel_data[5][103] = 4'b0111; // x=103, y=5
        pixel_data[5][104] = 4'b0111; // x=104, y=5
        pixel_data[5][105] = 4'b0111; // x=105, y=5
        pixel_data[5][106] = 4'b0111; // x=106, y=5
        pixel_data[5][107] = 4'b0111; // x=107, y=5
        pixel_data[5][108] = 4'b0111; // x=108, y=5
        pixel_data[5][109] = 4'b0111; // x=109, y=5
        pixel_data[5][110] = 4'b0111; // x=110, y=5
        pixel_data[5][111] = 4'b0111; // x=111, y=5
        pixel_data[5][112] = 4'b0111; // x=112, y=5
        pixel_data[5][113] = 4'b0111; // x=113, y=5
        pixel_data[5][114] = 4'b0111; // x=114, y=5
        pixel_data[5][115] = 4'b0111; // x=115, y=5
        pixel_data[5][116] = 4'b0111; // x=116, y=5
        pixel_data[5][117] = 4'b0111; // x=117, y=5
        pixel_data[5][118] = 4'b0111; // x=118, y=5
        pixel_data[5][119] = 4'b0111; // x=119, y=5
        pixel_data[5][120] = 4'b0111; // x=120, y=5
        pixel_data[5][121] = 4'b0111; // x=121, y=5
        pixel_data[5][122] = 4'b0111; // x=122, y=5
        pixel_data[5][123] = 4'b0111; // x=123, y=5
        pixel_data[5][124] = 4'b0111; // x=124, y=5
        pixel_data[5][125] = 4'b0111; // x=125, y=5
        pixel_data[5][126] = 4'b0111; // x=126, y=5
        pixel_data[5][127] = 4'b0111; // x=127, y=5
        pixel_data[5][128] = 4'b0111; // x=128, y=5
        pixel_data[5][129] = 4'b0111; // x=129, y=5
        pixel_data[5][130] = 4'b0111; // x=130, y=5
        pixel_data[5][131] = 4'b0111; // x=131, y=5
        pixel_data[5][132] = 4'b0111; // x=132, y=5
        pixel_data[5][133] = 4'b0111; // x=133, y=5
        pixel_data[5][134] = 4'b0111; // x=134, y=5
        pixel_data[5][135] = 4'b0111; // x=135, y=5
        pixel_data[5][136] = 4'b0111; // x=136, y=5
        pixel_data[5][137] = 4'b0111; // x=137, y=5
        pixel_data[5][138] = 4'b0111; // x=138, y=5
        pixel_data[5][139] = 4'b0111; // x=139, y=5
        pixel_data[5][140] = 4'b0111; // x=140, y=5
        pixel_data[5][141] = 4'b0111; // x=141, y=5
        pixel_data[5][142] = 4'b0111; // x=142, y=5
        pixel_data[5][143] = 4'b0111; // x=143, y=5
        pixel_data[5][144] = 4'b0111; // x=144, y=5
        pixel_data[5][145] = 4'b0111; // x=145, y=5
        pixel_data[5][146] = 4'b0111; // x=146, y=5
        pixel_data[5][147] = 4'b0111; // x=147, y=5
        pixel_data[5][148] = 4'b0111; // x=148, y=5
        pixel_data[5][149] = 4'b0111; // x=149, y=5
        pixel_data[5][150] = 4'b0111; // x=150, y=5
        pixel_data[5][151] = 4'b0111; // x=151, y=5
        pixel_data[5][152] = 4'b0111; // x=152, y=5
        pixel_data[5][153] = 4'b0111; // x=153, y=5
        pixel_data[5][154] = 4'b0111; // x=154, y=5
        pixel_data[5][155] = 4'b0111; // x=155, y=5
        pixel_data[5][156] = 4'b0111; // x=156, y=5
        pixel_data[5][157] = 4'b0111; // x=157, y=5
        pixel_data[5][158] = 4'b0111; // x=158, y=5
        pixel_data[5][159] = 4'b0111; // x=159, y=5
        pixel_data[5][160] = 4'b0111; // x=160, y=5
        pixel_data[5][161] = 4'b0111; // x=161, y=5
        pixel_data[5][162] = 4'b0111; // x=162, y=5
        pixel_data[5][163] = 4'b0111; // x=163, y=5
        pixel_data[5][164] = 4'b0111; // x=164, y=5
        pixel_data[5][165] = 4'b0111; // x=165, y=5
        pixel_data[5][166] = 4'b0111; // x=166, y=5
        pixel_data[5][167] = 4'b0111; // x=167, y=5
        pixel_data[5][168] = 4'b0111; // x=168, y=5
        pixel_data[5][169] = 4'b0111; // x=169, y=5
        pixel_data[5][170] = 4'b0111; // x=170, y=5
        pixel_data[5][171] = 4'b0111; // x=171, y=5
        pixel_data[5][172] = 4'b0111; // x=172, y=5
        pixel_data[5][173] = 4'b0111; // x=173, y=5
        pixel_data[5][174] = 4'b0111; // x=174, y=5
        pixel_data[5][175] = 4'b0111; // x=175, y=5
        pixel_data[5][176] = 4'b0111; // x=176, y=5
        pixel_data[5][177] = 4'b0111; // x=177, y=5
        pixel_data[5][178] = 4'b0111; // x=178, y=5
        pixel_data[5][179] = 4'b0111; // x=179, y=5
        pixel_data[6][0] = 4'b0111; // x=0, y=6
        pixel_data[6][1] = 4'b0111; // x=1, y=6
        pixel_data[6][2] = 4'b0111; // x=2, y=6
        pixel_data[6][3] = 4'b0111; // x=3, y=6
        pixel_data[6][4] = 4'b0111; // x=4, y=6
        pixel_data[6][5] = 4'b0111; // x=5, y=6
        pixel_data[6][6] = 4'b0111; // x=6, y=6
        pixel_data[6][7] = 4'b0111; // x=7, y=6
        pixel_data[6][8] = 4'b0111; // x=8, y=6
        pixel_data[6][9] = 4'b0111; // x=9, y=6
        pixel_data[6][10] = 4'b0111; // x=10, y=6
        pixel_data[6][11] = 4'b0111; // x=11, y=6
        pixel_data[6][12] = 4'b0111; // x=12, y=6
        pixel_data[6][13] = 4'b0111; // x=13, y=6
        pixel_data[6][14] = 4'b0111; // x=14, y=6
        pixel_data[6][15] = 4'b0111; // x=15, y=6
        pixel_data[6][16] = 4'b0111; // x=16, y=6
        pixel_data[6][17] = 4'b0111; // x=17, y=6
        pixel_data[6][18] = 4'b0111; // x=18, y=6
        pixel_data[6][19] = 4'b0111; // x=19, y=6
        pixel_data[6][20] = 4'b0111; // x=20, y=6
        pixel_data[6][21] = 4'b0111; // x=21, y=6
        pixel_data[6][22] = 4'b0111; // x=22, y=6
        pixel_data[6][23] = 4'b0111; // x=23, y=6
        pixel_data[6][24] = 4'b0111; // x=24, y=6
        pixel_data[6][25] = 4'b0111; // x=25, y=6
        pixel_data[6][26] = 4'b0111; // x=26, y=6
        pixel_data[6][27] = 4'b0111; // x=27, y=6
        pixel_data[6][28] = 4'b0111; // x=28, y=6
        pixel_data[6][29] = 4'b0111; // x=29, y=6
        pixel_data[6][30] = 4'b0111; // x=30, y=6
        pixel_data[6][31] = 4'b0111; // x=31, y=6
        pixel_data[6][32] = 4'b0111; // x=32, y=6
        pixel_data[6][33] = 4'b0111; // x=33, y=6
        pixel_data[6][34] = 4'b0111; // x=34, y=6
        pixel_data[6][35] = 4'b0111; // x=35, y=6
        pixel_data[6][36] = 4'b0111; // x=36, y=6
        pixel_data[6][37] = 4'b0111; // x=37, y=6
        pixel_data[6][38] = 4'b0111; // x=38, y=6
        pixel_data[6][39] = 4'b0111; // x=39, y=6
        pixel_data[6][40] = 4'b0111; // x=40, y=6
        pixel_data[6][41] = 4'b0111; // x=41, y=6
        pixel_data[6][42] = 4'b0111; // x=42, y=6
        pixel_data[6][43] = 4'b0111; // x=43, y=6
        pixel_data[6][44] = 4'b0111; // x=44, y=6
        pixel_data[6][45] = 4'b0111; // x=45, y=6
        pixel_data[6][46] = 4'b0111; // x=46, y=6
        pixel_data[6][47] = 4'b0111; // x=47, y=6
        pixel_data[6][48] = 4'b0111; // x=48, y=6
        pixel_data[6][49] = 4'b0111; // x=49, y=6
        pixel_data[6][50] = 4'b0111; // x=50, y=6
        pixel_data[6][51] = 4'b0111; // x=51, y=6
        pixel_data[6][52] = 4'b0111; // x=52, y=6
        pixel_data[6][53] = 4'b0111; // x=53, y=6
        pixel_data[6][54] = 4'b0111; // x=54, y=6
        pixel_data[6][55] = 4'b0111; // x=55, y=6
        pixel_data[6][56] = 4'b0111; // x=56, y=6
        pixel_data[6][57] = 4'b0111; // x=57, y=6
        pixel_data[6][58] = 4'b0111; // x=58, y=6
        pixel_data[6][59] = 4'b0111; // x=59, y=6
        pixel_data[6][60] = 4'b0111; // x=60, y=6
        pixel_data[6][61] = 4'b0111; // x=61, y=6
        pixel_data[6][62] = 4'b0111; // x=62, y=6
        pixel_data[6][63] = 4'b0111; // x=63, y=6
        pixel_data[6][64] = 4'b0111; // x=64, y=6
        pixel_data[6][65] = 4'b0111; // x=65, y=6
        pixel_data[6][66] = 4'b0111; // x=66, y=6
        pixel_data[6][67] = 4'b0111; // x=67, y=6
        pixel_data[6][68] = 4'b0111; // x=68, y=6
        pixel_data[6][69] = 4'b0111; // x=69, y=6
        pixel_data[6][70] = 4'b0111; // x=70, y=6
        pixel_data[6][71] = 4'b0111; // x=71, y=6
        pixel_data[6][72] = 4'b0111; // x=72, y=6
        pixel_data[6][73] = 4'b0111; // x=73, y=6
        pixel_data[6][74] = 4'b0111; // x=74, y=6
        pixel_data[6][75] = 4'b0111; // x=75, y=6
        pixel_data[6][76] = 4'b0111; // x=76, y=6
        pixel_data[6][77] = 4'b0111; // x=77, y=6
        pixel_data[6][78] = 4'b0111; // x=78, y=6
        pixel_data[6][79] = 4'b0111; // x=79, y=6
        pixel_data[6][80] = 4'b0111; // x=80, y=6
        pixel_data[6][81] = 4'b0111; // x=81, y=6
        pixel_data[6][82] = 4'b0111; // x=82, y=6
        pixel_data[6][83] = 4'b0111; // x=83, y=6
        pixel_data[6][84] = 4'b0111; // x=84, y=6
        pixel_data[6][85] = 4'b0111; // x=85, y=6
        pixel_data[6][86] = 4'b0111; // x=86, y=6
        pixel_data[6][87] = 4'b0111; // x=87, y=6
        pixel_data[6][88] = 4'b0111; // x=88, y=6
        pixel_data[6][89] = 4'b0111; // x=89, y=6
        pixel_data[6][90] = 4'b0111; // x=90, y=6
        pixel_data[6][91] = 4'b0111; // x=91, y=6
        pixel_data[6][92] = 4'b0111; // x=92, y=6
        pixel_data[6][93] = 4'b0111; // x=93, y=6
        pixel_data[6][94] = 4'b0111; // x=94, y=6
        pixel_data[6][95] = 4'b0111; // x=95, y=6
        pixel_data[6][96] = 4'b0111; // x=96, y=6
        pixel_data[6][97] = 4'b0111; // x=97, y=6
        pixel_data[6][98] = 4'b0111; // x=98, y=6
        pixel_data[6][99] = 4'b0111; // x=99, y=6
        pixel_data[6][100] = 4'b0111; // x=100, y=6
        pixel_data[6][101] = 4'b0111; // x=101, y=6
        pixel_data[6][102] = 4'b0111; // x=102, y=6
        pixel_data[6][103] = 4'b0111; // x=103, y=6
        pixel_data[6][104] = 4'b0111; // x=104, y=6
        pixel_data[6][105] = 4'b0111; // x=105, y=6
        pixel_data[6][106] = 4'b0111; // x=106, y=6
        pixel_data[6][107] = 4'b0111; // x=107, y=6
        pixel_data[6][108] = 4'b0111; // x=108, y=6
        pixel_data[6][109] = 4'b0111; // x=109, y=6
        pixel_data[6][110] = 4'b0111; // x=110, y=6
        pixel_data[6][111] = 4'b0111; // x=111, y=6
        pixel_data[6][112] = 4'b0111; // x=112, y=6
        pixel_data[6][113] = 4'b0111; // x=113, y=6
        pixel_data[6][114] = 4'b0111; // x=114, y=6
        pixel_data[6][115] = 4'b0111; // x=115, y=6
        pixel_data[6][116] = 4'b0111; // x=116, y=6
        pixel_data[6][117] = 4'b0111; // x=117, y=6
        pixel_data[6][118] = 4'b0111; // x=118, y=6
        pixel_data[6][119] = 4'b0111; // x=119, y=6
        pixel_data[6][120] = 4'b0111; // x=120, y=6
        pixel_data[6][121] = 4'b0111; // x=121, y=6
        pixel_data[6][122] = 4'b0111; // x=122, y=6
        pixel_data[6][123] = 4'b0111; // x=123, y=6
        pixel_data[6][124] = 4'b0111; // x=124, y=6
        pixel_data[6][125] = 4'b0111; // x=125, y=6
        pixel_data[6][126] = 4'b0111; // x=126, y=6
        pixel_data[6][127] = 4'b0111; // x=127, y=6
        pixel_data[6][128] = 4'b0111; // x=128, y=6
        pixel_data[6][129] = 4'b0111; // x=129, y=6
        pixel_data[6][130] = 4'b0111; // x=130, y=6
        pixel_data[6][131] = 4'b0111; // x=131, y=6
        pixel_data[6][132] = 4'b0111; // x=132, y=6
        pixel_data[6][133] = 4'b0111; // x=133, y=6
        pixel_data[6][134] = 4'b0111; // x=134, y=6
        pixel_data[6][135] = 4'b0111; // x=135, y=6
        pixel_data[6][136] = 4'b0111; // x=136, y=6
        pixel_data[6][137] = 4'b0111; // x=137, y=6
        pixel_data[6][138] = 4'b0111; // x=138, y=6
        pixel_data[6][139] = 4'b0111; // x=139, y=6
        pixel_data[6][140] = 4'b0111; // x=140, y=6
        pixel_data[6][141] = 4'b0111; // x=141, y=6
        pixel_data[6][142] = 4'b0111; // x=142, y=6
        pixel_data[6][143] = 4'b0111; // x=143, y=6
        pixel_data[6][144] = 4'b0111; // x=144, y=6
        pixel_data[6][145] = 4'b0111; // x=145, y=6
        pixel_data[6][146] = 4'b0111; // x=146, y=6
        pixel_data[6][147] = 4'b0111; // x=147, y=6
        pixel_data[6][148] = 4'b0111; // x=148, y=6
        pixel_data[6][149] = 4'b0111; // x=149, y=6
        pixel_data[6][150] = 4'b0111; // x=150, y=6
        pixel_data[6][151] = 4'b0111; // x=151, y=6
        pixel_data[6][152] = 4'b0111; // x=152, y=6
        pixel_data[6][153] = 4'b0111; // x=153, y=6
        pixel_data[6][154] = 4'b0111; // x=154, y=6
        pixel_data[6][155] = 4'b0111; // x=155, y=6
        pixel_data[6][156] = 4'b0111; // x=156, y=6
        pixel_data[6][157] = 4'b0111; // x=157, y=6
        pixel_data[6][158] = 4'b0111; // x=158, y=6
        pixel_data[6][159] = 4'b0111; // x=159, y=6
        pixel_data[6][160] = 4'b0111; // x=160, y=6
        pixel_data[6][161] = 4'b0111; // x=161, y=6
        pixel_data[6][162] = 4'b0111; // x=162, y=6
        pixel_data[6][163] = 4'b0111; // x=163, y=6
        pixel_data[6][164] = 4'b0111; // x=164, y=6
        pixel_data[6][165] = 4'b0111; // x=165, y=6
        pixel_data[6][166] = 4'b0111; // x=166, y=6
        pixel_data[6][167] = 4'b0111; // x=167, y=6
        pixel_data[6][168] = 4'b0111; // x=168, y=6
        pixel_data[6][169] = 4'b0111; // x=169, y=6
        pixel_data[6][170] = 4'b0111; // x=170, y=6
        pixel_data[6][171] = 4'b0111; // x=171, y=6
        pixel_data[6][172] = 4'b0111; // x=172, y=6
        pixel_data[6][173] = 4'b0111; // x=173, y=6
        pixel_data[6][174] = 4'b0111; // x=174, y=6
        pixel_data[6][175] = 4'b0111; // x=175, y=6
        pixel_data[6][176] = 4'b0111; // x=176, y=6
        pixel_data[6][177] = 4'b0111; // x=177, y=6
        pixel_data[6][178] = 4'b0111; // x=178, y=6
        pixel_data[6][179] = 4'b0111; // x=179, y=6
        pixel_data[7][0] = 4'b0111; // x=0, y=7
        pixel_data[7][1] = 4'b0111; // x=1, y=7
        pixel_data[7][2] = 4'b0111; // x=2, y=7
        pixel_data[7][3] = 4'b0111; // x=3, y=7
        pixel_data[7][4] = 4'b0111; // x=4, y=7
        pixel_data[7][5] = 4'b0111; // x=5, y=7
        pixel_data[7][6] = 4'b0111; // x=6, y=7
        pixel_data[7][7] = 4'b0111; // x=7, y=7
        pixel_data[7][8] = 4'b0111; // x=8, y=7
        pixel_data[7][9] = 4'b0111; // x=9, y=7
        pixel_data[7][10] = 4'b0111; // x=10, y=7
        pixel_data[7][11] = 4'b0111; // x=11, y=7
        pixel_data[7][12] = 4'b0111; // x=12, y=7
        pixel_data[7][13] = 4'b0111; // x=13, y=7
        pixel_data[7][14] = 4'b0111; // x=14, y=7
        pixel_data[7][15] = 4'b0111; // x=15, y=7
        pixel_data[7][16] = 4'b0111; // x=16, y=7
        pixel_data[7][17] = 4'b0111; // x=17, y=7
        pixel_data[7][18] = 4'b0111; // x=18, y=7
        pixel_data[7][19] = 4'b0111; // x=19, y=7
        pixel_data[7][20] = 4'b0111; // x=20, y=7
        pixel_data[7][21] = 4'b0111; // x=21, y=7
        pixel_data[7][22] = 4'b0111; // x=22, y=7
        pixel_data[7][23] = 4'b0111; // x=23, y=7
        pixel_data[7][24] = 4'b0111; // x=24, y=7
        pixel_data[7][25] = 4'b0111; // x=25, y=7
        pixel_data[7][26] = 4'b0111; // x=26, y=7
        pixel_data[7][27] = 4'b0111; // x=27, y=7
        pixel_data[7][28] = 4'b0111; // x=28, y=7
        pixel_data[7][29] = 4'b0111; // x=29, y=7
        pixel_data[7][30] = 4'b0111; // x=30, y=7
        pixel_data[7][31] = 4'b0111; // x=31, y=7
        pixel_data[7][32] = 4'b0111; // x=32, y=7
        pixel_data[7][33] = 4'b0111; // x=33, y=7
        pixel_data[7][34] = 4'b0111; // x=34, y=7
        pixel_data[7][35] = 4'b0111; // x=35, y=7
        pixel_data[7][36] = 4'b0111; // x=36, y=7
        pixel_data[7][37] = 4'b0111; // x=37, y=7
        pixel_data[7][38] = 4'b0111; // x=38, y=7
        pixel_data[7][39] = 4'b0111; // x=39, y=7
        pixel_data[7][40] = 4'b0111; // x=40, y=7
        pixel_data[7][41] = 4'b0111; // x=41, y=7
        pixel_data[7][42] = 4'b0111; // x=42, y=7
        pixel_data[7][43] = 4'b0111; // x=43, y=7
        pixel_data[7][44] = 4'b0111; // x=44, y=7
        pixel_data[7][45] = 4'b0111; // x=45, y=7
        pixel_data[7][46] = 4'b0111; // x=46, y=7
        pixel_data[7][47] = 4'b0111; // x=47, y=7
        pixel_data[7][48] = 4'b0111; // x=48, y=7
        pixel_data[7][49] = 4'b0111; // x=49, y=7
        pixel_data[7][50] = 4'b0111; // x=50, y=7
        pixel_data[7][51] = 4'b0111; // x=51, y=7
        pixel_data[7][52] = 4'b0111; // x=52, y=7
        pixel_data[7][53] = 4'b0111; // x=53, y=7
        pixel_data[7][54] = 4'b0111; // x=54, y=7
        pixel_data[7][55] = 4'b0111; // x=55, y=7
        pixel_data[7][56] = 4'b0111; // x=56, y=7
        pixel_data[7][57] = 4'b0111; // x=57, y=7
        pixel_data[7][58] = 4'b0111; // x=58, y=7
        pixel_data[7][59] = 4'b0111; // x=59, y=7
        pixel_data[7][60] = 4'b0111; // x=60, y=7
        pixel_data[7][61] = 4'b0111; // x=61, y=7
        pixel_data[7][62] = 4'b0111; // x=62, y=7
        pixel_data[7][63] = 4'b0111; // x=63, y=7
        pixel_data[7][64] = 4'b0111; // x=64, y=7
        pixel_data[7][65] = 4'b0111; // x=65, y=7
        pixel_data[7][66] = 4'b0111; // x=66, y=7
        pixel_data[7][67] = 4'b0111; // x=67, y=7
        pixel_data[7][68] = 4'b0111; // x=68, y=7
        pixel_data[7][69] = 4'b0111; // x=69, y=7
        pixel_data[7][70] = 4'b0111; // x=70, y=7
        pixel_data[7][71] = 4'b0111; // x=71, y=7
        pixel_data[7][72] = 4'b0111; // x=72, y=7
        pixel_data[7][73] = 4'b0111; // x=73, y=7
        pixel_data[7][74] = 4'b0111; // x=74, y=7
        pixel_data[7][75] = 4'b0111; // x=75, y=7
        pixel_data[7][76] = 4'b0111; // x=76, y=7
        pixel_data[7][77] = 4'b0111; // x=77, y=7
        pixel_data[7][78] = 4'b0111; // x=78, y=7
        pixel_data[7][79] = 4'b0111; // x=79, y=7
        pixel_data[7][80] = 4'b0111; // x=80, y=7
        pixel_data[7][81] = 4'b0111; // x=81, y=7
        pixel_data[7][82] = 4'b0111; // x=82, y=7
        pixel_data[7][83] = 4'b0111; // x=83, y=7
        pixel_data[7][84] = 4'b0111; // x=84, y=7
        pixel_data[7][85] = 4'b0111; // x=85, y=7
        pixel_data[7][86] = 4'b0111; // x=86, y=7
        pixel_data[7][87] = 4'b0111; // x=87, y=7
        pixel_data[7][88] = 4'b0111; // x=88, y=7
        pixel_data[7][89] = 4'b0111; // x=89, y=7
        pixel_data[7][90] = 4'b0111; // x=90, y=7
        pixel_data[7][91] = 4'b0111; // x=91, y=7
        pixel_data[7][92] = 4'b0111; // x=92, y=7
        pixel_data[7][93] = 4'b0111; // x=93, y=7
        pixel_data[7][94] = 4'b0111; // x=94, y=7
        pixel_data[7][95] = 4'b0111; // x=95, y=7
        pixel_data[7][96] = 4'b0111; // x=96, y=7
        pixel_data[7][97] = 4'b0111; // x=97, y=7
        pixel_data[7][98] = 4'b0111; // x=98, y=7
        pixel_data[7][99] = 4'b0111; // x=99, y=7
        pixel_data[7][100] = 4'b0111; // x=100, y=7
        pixel_data[7][101] = 4'b0111; // x=101, y=7
        pixel_data[7][102] = 4'b0111; // x=102, y=7
        pixel_data[7][103] = 4'b0111; // x=103, y=7
        pixel_data[7][104] = 4'b0111; // x=104, y=7
        pixel_data[7][105] = 4'b0111; // x=105, y=7
        pixel_data[7][106] = 4'b0111; // x=106, y=7
        pixel_data[7][107] = 4'b0111; // x=107, y=7
        pixel_data[7][108] = 4'b0111; // x=108, y=7
        pixel_data[7][109] = 4'b0111; // x=109, y=7
        pixel_data[7][110] = 4'b0111; // x=110, y=7
        pixel_data[7][111] = 4'b0111; // x=111, y=7
        pixel_data[7][112] = 4'b0111; // x=112, y=7
        pixel_data[7][113] = 4'b0111; // x=113, y=7
        pixel_data[7][114] = 4'b0111; // x=114, y=7
        pixel_data[7][115] = 4'b0111; // x=115, y=7
        pixel_data[7][116] = 4'b0111; // x=116, y=7
        pixel_data[7][117] = 4'b0111; // x=117, y=7
        pixel_data[7][118] = 4'b0111; // x=118, y=7
        pixel_data[7][119] = 4'b0111; // x=119, y=7
        pixel_data[7][120] = 4'b0111; // x=120, y=7
        pixel_data[7][121] = 4'b0111; // x=121, y=7
        pixel_data[7][122] = 4'b0111; // x=122, y=7
        pixel_data[7][123] = 4'b0111; // x=123, y=7
        pixel_data[7][124] = 4'b0111; // x=124, y=7
        pixel_data[7][125] = 4'b0111; // x=125, y=7
        pixel_data[7][126] = 4'b0111; // x=126, y=7
        pixel_data[7][127] = 4'b0111; // x=127, y=7
        pixel_data[7][128] = 4'b0111; // x=128, y=7
        pixel_data[7][129] = 4'b0111; // x=129, y=7
        pixel_data[7][130] = 4'b0111; // x=130, y=7
        pixel_data[7][131] = 4'b0111; // x=131, y=7
        pixel_data[7][132] = 4'b0111; // x=132, y=7
        pixel_data[7][133] = 4'b0111; // x=133, y=7
        pixel_data[7][134] = 4'b0111; // x=134, y=7
        pixel_data[7][135] = 4'b0111; // x=135, y=7
        pixel_data[7][136] = 4'b0111; // x=136, y=7
        pixel_data[7][137] = 4'b0111; // x=137, y=7
        pixel_data[7][138] = 4'b0111; // x=138, y=7
        pixel_data[7][139] = 4'b0111; // x=139, y=7
        pixel_data[7][140] = 4'b0111; // x=140, y=7
        pixel_data[7][141] = 4'b0111; // x=141, y=7
        pixel_data[7][142] = 4'b0111; // x=142, y=7
        pixel_data[7][143] = 4'b0111; // x=143, y=7
        pixel_data[7][144] = 4'b0111; // x=144, y=7
        pixel_data[7][145] = 4'b0111; // x=145, y=7
        pixel_data[7][146] = 4'b0111; // x=146, y=7
        pixel_data[7][147] = 4'b0111; // x=147, y=7
        pixel_data[7][148] = 4'b0111; // x=148, y=7
        pixel_data[7][149] = 4'b0111; // x=149, y=7
        pixel_data[7][150] = 4'b0111; // x=150, y=7
        pixel_data[7][151] = 4'b0111; // x=151, y=7
        pixel_data[7][152] = 4'b0111; // x=152, y=7
        pixel_data[7][153] = 4'b0111; // x=153, y=7
        pixel_data[7][154] = 4'b0111; // x=154, y=7
        pixel_data[7][155] = 4'b0111; // x=155, y=7
        pixel_data[7][156] = 4'b0111; // x=156, y=7
        pixel_data[7][157] = 4'b0111; // x=157, y=7
        pixel_data[7][158] = 4'b0111; // x=158, y=7
        pixel_data[7][159] = 4'b0111; // x=159, y=7
        pixel_data[7][160] = 4'b0111; // x=160, y=7
        pixel_data[7][161] = 4'b0111; // x=161, y=7
        pixel_data[7][162] = 4'b0111; // x=162, y=7
        pixel_data[7][163] = 4'b0111; // x=163, y=7
        pixel_data[7][164] = 4'b0111; // x=164, y=7
        pixel_data[7][165] = 4'b0111; // x=165, y=7
        pixel_data[7][166] = 4'b0111; // x=166, y=7
        pixel_data[7][167] = 4'b0111; // x=167, y=7
        pixel_data[7][168] = 4'b0111; // x=168, y=7
        pixel_data[7][169] = 4'b0111; // x=169, y=7
        pixel_data[7][170] = 4'b0111; // x=170, y=7
        pixel_data[7][171] = 4'b0111; // x=171, y=7
        pixel_data[7][172] = 4'b0111; // x=172, y=7
        pixel_data[7][173] = 4'b0111; // x=173, y=7
        pixel_data[7][174] = 4'b0111; // x=174, y=7
        pixel_data[7][175] = 4'b0111; // x=175, y=7
        pixel_data[7][176] = 4'b0111; // x=176, y=7
        pixel_data[7][177] = 4'b0111; // x=177, y=7
        pixel_data[7][178] = 4'b0111; // x=178, y=7
        pixel_data[7][179] = 4'b0111; // x=179, y=7
        pixel_data[8][0] = 4'b0111; // x=0, y=8
        pixel_data[8][1] = 4'b0111; // x=1, y=8
        pixel_data[8][2] = 4'b0111; // x=2, y=8
        pixel_data[8][3] = 4'b0111; // x=3, y=8
        pixel_data[8][4] = 4'b0111; // x=4, y=8
        pixel_data[8][5] = 4'b0111; // x=5, y=8
        pixel_data[8][6] = 4'b0111; // x=6, y=8
        pixel_data[8][7] = 4'b0111; // x=7, y=8
        pixel_data[8][8] = 4'b0111; // x=8, y=8
        pixel_data[8][9] = 4'b0111; // x=9, y=8
        pixel_data[8][10] = 4'b0111; // x=10, y=8
        pixel_data[8][11] = 4'b0111; // x=11, y=8
        pixel_data[8][12] = 4'b0111; // x=12, y=8
        pixel_data[8][13] = 4'b0111; // x=13, y=8
        pixel_data[8][14] = 4'b0111; // x=14, y=8
        pixel_data[8][15] = 4'b0111; // x=15, y=8
        pixel_data[8][16] = 4'b0111; // x=16, y=8
        pixel_data[8][17] = 4'b0111; // x=17, y=8
        pixel_data[8][18] = 4'b0111; // x=18, y=8
        pixel_data[8][19] = 4'b0111; // x=19, y=8
        pixel_data[8][20] = 4'b0111; // x=20, y=8
        pixel_data[8][21] = 4'b0111; // x=21, y=8
        pixel_data[8][22] = 4'b0111; // x=22, y=8
        pixel_data[8][23] = 4'b0111; // x=23, y=8
        pixel_data[8][24] = 4'b0111; // x=24, y=8
        pixel_data[8][25] = 4'b0111; // x=25, y=8
        pixel_data[8][26] = 4'b0111; // x=26, y=8
        pixel_data[8][27] = 4'b0111; // x=27, y=8
        pixel_data[8][28] = 4'b0111; // x=28, y=8
        pixel_data[8][29] = 4'b0111; // x=29, y=8
        pixel_data[8][30] = 4'b0111; // x=30, y=8
        pixel_data[8][31] = 4'b0111; // x=31, y=8
        pixel_data[8][32] = 4'b0111; // x=32, y=8
        pixel_data[8][33] = 4'b0111; // x=33, y=8
        pixel_data[8][34] = 4'b0111; // x=34, y=8
        pixel_data[8][35] = 4'b0111; // x=35, y=8
        pixel_data[8][36] = 4'b0111; // x=36, y=8
        pixel_data[8][37] = 4'b0111; // x=37, y=8
        pixel_data[8][38] = 4'b0111; // x=38, y=8
        pixel_data[8][39] = 4'b0111; // x=39, y=8
        pixel_data[8][40] = 4'b0111; // x=40, y=8
        pixel_data[8][41] = 4'b0111; // x=41, y=8
        pixel_data[8][42] = 4'b0111; // x=42, y=8
        pixel_data[8][43] = 4'b0111; // x=43, y=8
        pixel_data[8][44] = 4'b0111; // x=44, y=8
        pixel_data[8][45] = 4'b0111; // x=45, y=8
        pixel_data[8][46] = 4'b0111; // x=46, y=8
        pixel_data[8][47] = 4'b0111; // x=47, y=8
        pixel_data[8][48] = 4'b0111; // x=48, y=8
        pixel_data[8][49] = 4'b0111; // x=49, y=8
        pixel_data[8][50] = 4'b0111; // x=50, y=8
        pixel_data[8][51] = 4'b0111; // x=51, y=8
        pixel_data[8][52] = 4'b0111; // x=52, y=8
        pixel_data[8][53] = 4'b0111; // x=53, y=8
        pixel_data[8][54] = 4'b0111; // x=54, y=8
        pixel_data[8][55] = 4'b0111; // x=55, y=8
        pixel_data[8][56] = 4'b0111; // x=56, y=8
        pixel_data[8][57] = 4'b0111; // x=57, y=8
        pixel_data[8][58] = 4'b0111; // x=58, y=8
        pixel_data[8][59] = 4'b0111; // x=59, y=8
        pixel_data[8][60] = 4'b0111; // x=60, y=8
        pixel_data[8][61] = 4'b0111; // x=61, y=8
        pixel_data[8][62] = 4'b0111; // x=62, y=8
        pixel_data[8][63] = 4'b0111; // x=63, y=8
        pixel_data[8][64] = 4'b0111; // x=64, y=8
        pixel_data[8][65] = 4'b0111; // x=65, y=8
        pixel_data[8][66] = 4'b0111; // x=66, y=8
        pixel_data[8][67] = 4'b0111; // x=67, y=8
        pixel_data[8][68] = 4'b0111; // x=68, y=8
        pixel_data[8][69] = 4'b0111; // x=69, y=8
        pixel_data[8][70] = 4'b0111; // x=70, y=8
        pixel_data[8][71] = 4'b0111; // x=71, y=8
        pixel_data[8][72] = 4'b0111; // x=72, y=8
        pixel_data[8][73] = 4'b0111; // x=73, y=8
        pixel_data[8][74] = 4'b0111; // x=74, y=8
        pixel_data[8][75] = 4'b0111; // x=75, y=8
        pixel_data[8][76] = 4'b0111; // x=76, y=8
        pixel_data[8][77] = 4'b0111; // x=77, y=8
        pixel_data[8][78] = 4'b0111; // x=78, y=8
        pixel_data[8][79] = 4'b0111; // x=79, y=8
        pixel_data[8][80] = 4'b0111; // x=80, y=8
        pixel_data[8][81] = 4'b0111; // x=81, y=8
        pixel_data[8][82] = 4'b0111; // x=82, y=8
        pixel_data[8][83] = 4'b0111; // x=83, y=8
        pixel_data[8][84] = 4'b0111; // x=84, y=8
        pixel_data[8][85] = 4'b0111; // x=85, y=8
        pixel_data[8][86] = 4'b0111; // x=86, y=8
        pixel_data[8][87] = 4'b0111; // x=87, y=8
        pixel_data[8][88] = 4'b0111; // x=88, y=8
        pixel_data[8][89] = 4'b0111; // x=89, y=8
        pixel_data[8][90] = 4'b0111; // x=90, y=8
        pixel_data[8][91] = 4'b0111; // x=91, y=8
        pixel_data[8][92] = 4'b0111; // x=92, y=8
        pixel_data[8][93] = 4'b0111; // x=93, y=8
        pixel_data[8][94] = 4'b0111; // x=94, y=8
        pixel_data[8][95] = 4'b0111; // x=95, y=8
        pixel_data[8][96] = 4'b0111; // x=96, y=8
        pixel_data[8][97] = 4'b0111; // x=97, y=8
        pixel_data[8][98] = 4'b0111; // x=98, y=8
        pixel_data[8][99] = 4'b0111; // x=99, y=8
        pixel_data[8][100] = 4'b0111; // x=100, y=8
        pixel_data[8][101] = 4'b0111; // x=101, y=8
        pixel_data[8][102] = 4'b0111; // x=102, y=8
        pixel_data[8][103] = 4'b0111; // x=103, y=8
        pixel_data[8][104] = 4'b0111; // x=104, y=8
        pixel_data[8][105] = 4'b0111; // x=105, y=8
        pixel_data[8][106] = 4'b0111; // x=106, y=8
        pixel_data[8][107] = 4'b0111; // x=107, y=8
        pixel_data[8][108] = 4'b0111; // x=108, y=8
        pixel_data[8][109] = 4'b0111; // x=109, y=8
        pixel_data[8][110] = 4'b0111; // x=110, y=8
        pixel_data[8][111] = 4'b0111; // x=111, y=8
        pixel_data[8][112] = 4'b0111; // x=112, y=8
        pixel_data[8][113] = 4'b0111; // x=113, y=8
        pixel_data[8][114] = 4'b0111; // x=114, y=8
        pixel_data[8][115] = 4'b0111; // x=115, y=8
        pixel_data[8][116] = 4'b0111; // x=116, y=8
        pixel_data[8][117] = 4'b0111; // x=117, y=8
        pixel_data[8][118] = 4'b0111; // x=118, y=8
        pixel_data[8][119] = 4'b0111; // x=119, y=8
        pixel_data[8][120] = 4'b0111; // x=120, y=8
        pixel_data[8][121] = 4'b0111; // x=121, y=8
        pixel_data[8][122] = 4'b0111; // x=122, y=8
        pixel_data[8][123] = 4'b0111; // x=123, y=8
        pixel_data[8][124] = 4'b0111; // x=124, y=8
        pixel_data[8][125] = 4'b0111; // x=125, y=8
        pixel_data[8][126] = 4'b0111; // x=126, y=8
        pixel_data[8][127] = 4'b0111; // x=127, y=8
        pixel_data[8][128] = 4'b0111; // x=128, y=8
        pixel_data[8][129] = 4'b0111; // x=129, y=8
        pixel_data[8][130] = 4'b0111; // x=130, y=8
        pixel_data[8][131] = 4'b0111; // x=131, y=8
        pixel_data[8][132] = 4'b0111; // x=132, y=8
        pixel_data[8][133] = 4'b0111; // x=133, y=8
        pixel_data[8][134] = 4'b0111; // x=134, y=8
        pixel_data[8][135] = 4'b0111; // x=135, y=8
        pixel_data[8][136] = 4'b0111; // x=136, y=8
        pixel_data[8][137] = 4'b0111; // x=137, y=8
        pixel_data[8][138] = 4'b0111; // x=138, y=8
        pixel_data[8][139] = 4'b0111; // x=139, y=8
        pixel_data[8][140] = 4'b0111; // x=140, y=8
        pixel_data[8][141] = 4'b0111; // x=141, y=8
        pixel_data[8][142] = 4'b0111; // x=142, y=8
        pixel_data[8][143] = 4'b0111; // x=143, y=8
        pixel_data[8][144] = 4'b0111; // x=144, y=8
        pixel_data[8][145] = 4'b0111; // x=145, y=8
        pixel_data[8][146] = 4'b0111; // x=146, y=8
        pixel_data[8][147] = 4'b0111; // x=147, y=8
        pixel_data[8][148] = 4'b0111; // x=148, y=8
        pixel_data[8][149] = 4'b0111; // x=149, y=8
        pixel_data[8][150] = 4'b0111; // x=150, y=8
        pixel_data[8][151] = 4'b0111; // x=151, y=8
        pixel_data[8][152] = 4'b0111; // x=152, y=8
        pixel_data[8][153] = 4'b0111; // x=153, y=8
        pixel_data[8][154] = 4'b0111; // x=154, y=8
        pixel_data[8][155] = 4'b0111; // x=155, y=8
        pixel_data[8][156] = 4'b0111; // x=156, y=8
        pixel_data[8][157] = 4'b0111; // x=157, y=8
        pixel_data[8][158] = 4'b0111; // x=158, y=8
        pixel_data[8][159] = 4'b0111; // x=159, y=8
        pixel_data[8][160] = 4'b0111; // x=160, y=8
        pixel_data[8][161] = 4'b0111; // x=161, y=8
        pixel_data[8][162] = 4'b0111; // x=162, y=8
        pixel_data[8][163] = 4'b0111; // x=163, y=8
        pixel_data[8][164] = 4'b0111; // x=164, y=8
        pixel_data[8][165] = 4'b0111; // x=165, y=8
        pixel_data[8][166] = 4'b0111; // x=166, y=8
        pixel_data[8][167] = 4'b0111; // x=167, y=8
        pixel_data[8][168] = 4'b0111; // x=168, y=8
        pixel_data[8][169] = 4'b0111; // x=169, y=8
        pixel_data[8][170] = 4'b0111; // x=170, y=8
        pixel_data[8][171] = 4'b0111; // x=171, y=8
        pixel_data[8][172] = 4'b0111; // x=172, y=8
        pixel_data[8][173] = 4'b0111; // x=173, y=8
        pixel_data[8][174] = 4'b0111; // x=174, y=8
        pixel_data[8][175] = 4'b0111; // x=175, y=8
        pixel_data[8][176] = 4'b0111; // x=176, y=8
        pixel_data[8][177] = 4'b0111; // x=177, y=8
        pixel_data[8][178] = 4'b0111; // x=178, y=8
        pixel_data[8][179] = 4'b0111; // x=179, y=8
        pixel_data[9][0] = 4'b0111; // x=0, y=9
        pixel_data[9][1] = 4'b0111; // x=1, y=9
        pixel_data[9][2] = 4'b0111; // x=2, y=9
        pixel_data[9][3] = 4'b0111; // x=3, y=9
        pixel_data[9][4] = 4'b0111; // x=4, y=9
        pixel_data[9][5] = 4'b0111; // x=5, y=9
        pixel_data[9][6] = 4'b0111; // x=6, y=9
        pixel_data[9][7] = 4'b0111; // x=7, y=9
        pixel_data[9][8] = 4'b0111; // x=8, y=9
        pixel_data[9][9] = 4'b0111; // x=9, y=9
        pixel_data[9][10] = 4'b0111; // x=10, y=9
        pixel_data[9][11] = 4'b0111; // x=11, y=9
        pixel_data[9][12] = 4'b0111; // x=12, y=9
        pixel_data[9][13] = 4'b0111; // x=13, y=9
        pixel_data[9][14] = 4'b0111; // x=14, y=9
        pixel_data[9][15] = 4'b0111; // x=15, y=9
        pixel_data[9][16] = 4'b0111; // x=16, y=9
        pixel_data[9][17] = 4'b0111; // x=17, y=9
        pixel_data[9][18] = 4'b0111; // x=18, y=9
        pixel_data[9][19] = 4'b0111; // x=19, y=9
        pixel_data[9][20] = 4'b0111; // x=20, y=9
        pixel_data[9][21] = 4'b0111; // x=21, y=9
        pixel_data[9][22] = 4'b0111; // x=22, y=9
        pixel_data[9][23] = 4'b0111; // x=23, y=9
        pixel_data[9][24] = 4'b0111; // x=24, y=9
        pixel_data[9][25] = 4'b0111; // x=25, y=9
        pixel_data[9][26] = 4'b0111; // x=26, y=9
        pixel_data[9][27] = 4'b0111; // x=27, y=9
        pixel_data[9][28] = 4'b0111; // x=28, y=9
        pixel_data[9][29] = 4'b0111; // x=29, y=9
        pixel_data[9][30] = 4'b0111; // x=30, y=9
        pixel_data[9][31] = 4'b0111; // x=31, y=9
        pixel_data[9][32] = 4'b0111; // x=32, y=9
        pixel_data[9][33] = 4'b0111; // x=33, y=9
        pixel_data[9][34] = 4'b0111; // x=34, y=9
        pixel_data[9][35] = 4'b0111; // x=35, y=9
        pixel_data[9][36] = 4'b0111; // x=36, y=9
        pixel_data[9][37] = 4'b0111; // x=37, y=9
        pixel_data[9][38] = 4'b0111; // x=38, y=9
        pixel_data[9][39] = 4'b0111; // x=39, y=9
        pixel_data[9][40] = 4'b0111; // x=40, y=9
        pixel_data[9][41] = 4'b0111; // x=41, y=9
        pixel_data[9][42] = 4'b0111; // x=42, y=9
        pixel_data[9][43] = 4'b0111; // x=43, y=9
        pixel_data[9][44] = 4'b0111; // x=44, y=9
        pixel_data[9][45] = 4'b0111; // x=45, y=9
        pixel_data[9][46] = 4'b0111; // x=46, y=9
        pixel_data[9][47] = 4'b0111; // x=47, y=9
        pixel_data[9][48] = 4'b0111; // x=48, y=9
        pixel_data[9][49] = 4'b0111; // x=49, y=9
        pixel_data[9][50] = 4'b0111; // x=50, y=9
        pixel_data[9][51] = 4'b0111; // x=51, y=9
        pixel_data[9][52] = 4'b0111; // x=52, y=9
        pixel_data[9][53] = 4'b0111; // x=53, y=9
        pixel_data[9][54] = 4'b0111; // x=54, y=9
        pixel_data[9][55] = 4'b0111; // x=55, y=9
        pixel_data[9][56] = 4'b0111; // x=56, y=9
        pixel_data[9][57] = 4'b0111; // x=57, y=9
        pixel_data[9][58] = 4'b0111; // x=58, y=9
        pixel_data[9][59] = 4'b0111; // x=59, y=9
        pixel_data[9][60] = 4'b0111; // x=60, y=9
        pixel_data[9][61] = 4'b0111; // x=61, y=9
        pixel_data[9][62] = 4'b0111; // x=62, y=9
        pixel_data[9][63] = 4'b0111; // x=63, y=9
        pixel_data[9][64] = 4'b0111; // x=64, y=9
        pixel_data[9][65] = 4'b0111; // x=65, y=9
        pixel_data[9][66] = 4'b0111; // x=66, y=9
        pixel_data[9][67] = 4'b0111; // x=67, y=9
        pixel_data[9][68] = 4'b0111; // x=68, y=9
        pixel_data[9][69] = 4'b0111; // x=69, y=9
        pixel_data[9][70] = 4'b0111; // x=70, y=9
        pixel_data[9][71] = 4'b0111; // x=71, y=9
        pixel_data[9][72] = 4'b0111; // x=72, y=9
        pixel_data[9][73] = 4'b0111; // x=73, y=9
        pixel_data[9][74] = 4'b0111; // x=74, y=9
        pixel_data[9][75] = 4'b0111; // x=75, y=9
        pixel_data[9][76] = 4'b0111; // x=76, y=9
        pixel_data[9][77] = 4'b0111; // x=77, y=9
        pixel_data[9][78] = 4'b0111; // x=78, y=9
        pixel_data[9][79] = 4'b0111; // x=79, y=9
        pixel_data[9][80] = 4'b0111; // x=80, y=9
        pixel_data[9][81] = 4'b0111; // x=81, y=9
        pixel_data[9][82] = 4'b0111; // x=82, y=9
        pixel_data[9][83] = 4'b0111; // x=83, y=9
        pixel_data[9][84] = 4'b0111; // x=84, y=9
        pixel_data[9][85] = 4'b0111; // x=85, y=9
        pixel_data[9][86] = 4'b0111; // x=86, y=9
        pixel_data[9][87] = 4'b0111; // x=87, y=9
        pixel_data[9][88] = 4'b0111; // x=88, y=9
        pixel_data[9][89] = 4'b0111; // x=89, y=9
        pixel_data[9][90] = 4'b0111; // x=90, y=9
        pixel_data[9][91] = 4'b0111; // x=91, y=9
        pixel_data[9][92] = 4'b0111; // x=92, y=9
        pixel_data[9][93] = 4'b0111; // x=93, y=9
        pixel_data[9][94] = 4'b0111; // x=94, y=9
        pixel_data[9][95] = 4'b0111; // x=95, y=9
        pixel_data[9][96] = 4'b0111; // x=96, y=9
        pixel_data[9][97] = 4'b0111; // x=97, y=9
        pixel_data[9][98] = 4'b0111; // x=98, y=9
        pixel_data[9][99] = 4'b0111; // x=99, y=9
        pixel_data[9][100] = 4'b0111; // x=100, y=9
        pixel_data[9][101] = 4'b0111; // x=101, y=9
        pixel_data[9][102] = 4'b0111; // x=102, y=9
        pixel_data[9][103] = 4'b0111; // x=103, y=9
        pixel_data[9][104] = 4'b0111; // x=104, y=9
        pixel_data[9][105] = 4'b0111; // x=105, y=9
        pixel_data[9][106] = 4'b0111; // x=106, y=9
        pixel_data[9][107] = 4'b0111; // x=107, y=9
        pixel_data[9][108] = 4'b0111; // x=108, y=9
        pixel_data[9][109] = 4'b0111; // x=109, y=9
        pixel_data[9][110] = 4'b0111; // x=110, y=9
        pixel_data[9][111] = 4'b0111; // x=111, y=9
        pixel_data[9][112] = 4'b0111; // x=112, y=9
        pixel_data[9][113] = 4'b0111; // x=113, y=9
        pixel_data[9][114] = 4'b0111; // x=114, y=9
        pixel_data[9][115] = 4'b0111; // x=115, y=9
        pixel_data[9][116] = 4'b0111; // x=116, y=9
        pixel_data[9][117] = 4'b0111; // x=117, y=9
        pixel_data[9][118] = 4'b0111; // x=118, y=9
        pixel_data[9][119] = 4'b0111; // x=119, y=9
        pixel_data[9][120] = 4'b0111; // x=120, y=9
        pixel_data[9][121] = 4'b0111; // x=121, y=9
        pixel_data[9][122] = 4'b0111; // x=122, y=9
        pixel_data[9][123] = 4'b0111; // x=123, y=9
        pixel_data[9][124] = 4'b0111; // x=124, y=9
        pixel_data[9][125] = 4'b0111; // x=125, y=9
        pixel_data[9][126] = 4'b0111; // x=126, y=9
        pixel_data[9][127] = 4'b0111; // x=127, y=9
        pixel_data[9][128] = 4'b0111; // x=128, y=9
        pixel_data[9][129] = 4'b0111; // x=129, y=9
        pixel_data[9][130] = 4'b0111; // x=130, y=9
        pixel_data[9][131] = 4'b0111; // x=131, y=9
        pixel_data[9][132] = 4'b0111; // x=132, y=9
        pixel_data[9][133] = 4'b0111; // x=133, y=9
        pixel_data[9][134] = 4'b0111; // x=134, y=9
        pixel_data[9][135] = 4'b0111; // x=135, y=9
        pixel_data[9][136] = 4'b0111; // x=136, y=9
        pixel_data[9][137] = 4'b0111; // x=137, y=9
        pixel_data[9][138] = 4'b0111; // x=138, y=9
        pixel_data[9][139] = 4'b0111; // x=139, y=9
        pixel_data[9][140] = 4'b0111; // x=140, y=9
        pixel_data[9][141] = 4'b0111; // x=141, y=9
        pixel_data[9][142] = 4'b0111; // x=142, y=9
        pixel_data[9][143] = 4'b0111; // x=143, y=9
        pixel_data[9][144] = 4'b0111; // x=144, y=9
        pixel_data[9][145] = 4'b0111; // x=145, y=9
        pixel_data[9][146] = 4'b0111; // x=146, y=9
        pixel_data[9][147] = 4'b0111; // x=147, y=9
        pixel_data[9][148] = 4'b0111; // x=148, y=9
        pixel_data[9][149] = 4'b0111; // x=149, y=9
        pixel_data[9][150] = 4'b0111; // x=150, y=9
        pixel_data[9][151] = 4'b0111; // x=151, y=9
        pixel_data[9][152] = 4'b0111; // x=152, y=9
        pixel_data[9][153] = 4'b0111; // x=153, y=9
        pixel_data[9][154] = 4'b0111; // x=154, y=9
        pixel_data[9][155] = 4'b0111; // x=155, y=9
        pixel_data[9][156] = 4'b0111; // x=156, y=9
        pixel_data[9][157] = 4'b0111; // x=157, y=9
        pixel_data[9][158] = 4'b0111; // x=158, y=9
        pixel_data[9][159] = 4'b0111; // x=159, y=9
        pixel_data[9][160] = 4'b0111; // x=160, y=9
        pixel_data[9][161] = 4'b0111; // x=161, y=9
        pixel_data[9][162] = 4'b0111; // x=162, y=9
        pixel_data[9][163] = 4'b0111; // x=163, y=9
        pixel_data[9][164] = 4'b0111; // x=164, y=9
        pixel_data[9][165] = 4'b0111; // x=165, y=9
        pixel_data[9][166] = 4'b0111; // x=166, y=9
        pixel_data[9][167] = 4'b0111; // x=167, y=9
        pixel_data[9][168] = 4'b0111; // x=168, y=9
        pixel_data[9][169] = 4'b0111; // x=169, y=9
        pixel_data[9][170] = 4'b0111; // x=170, y=9
        pixel_data[9][171] = 4'b0111; // x=171, y=9
        pixel_data[9][172] = 4'b0111; // x=172, y=9
        pixel_data[9][173] = 4'b0111; // x=173, y=9
        pixel_data[9][174] = 4'b0111; // x=174, y=9
        pixel_data[9][175] = 4'b0111; // x=175, y=9
        pixel_data[9][176] = 4'b0111; // x=176, y=9
        pixel_data[9][177] = 4'b0111; // x=177, y=9
        pixel_data[9][178] = 4'b0111; // x=178, y=9
        pixel_data[9][179] = 4'b0111; // x=179, y=9
        pixel_data[10][0] = 4'b0111; // x=0, y=10
        pixel_data[10][1] = 4'b0111; // x=1, y=10
        pixel_data[10][2] = 4'b0111; // x=2, y=10
        pixel_data[10][3] = 4'b0111; // x=3, y=10
        pixel_data[10][4] = 4'b0111; // x=4, y=10
        pixel_data[10][5] = 4'b0111; // x=5, y=10
        pixel_data[10][6] = 4'b0111; // x=6, y=10
        pixel_data[10][7] = 4'b0111; // x=7, y=10
        pixel_data[10][8] = 4'b0111; // x=8, y=10
        pixel_data[10][9] = 4'b0111; // x=9, y=10
        pixel_data[10][10] = 4'b0111; // x=10, y=10
        pixel_data[10][11] = 4'b0111; // x=11, y=10
        pixel_data[10][12] = 4'b0111; // x=12, y=10
        pixel_data[10][13] = 4'b0111; // x=13, y=10
        pixel_data[10][14] = 4'b0111; // x=14, y=10
        pixel_data[10][15] = 4'b0111; // x=15, y=10
        pixel_data[10][16] = 4'b0111; // x=16, y=10
        pixel_data[10][17] = 4'b0111; // x=17, y=10
        pixel_data[10][18] = 4'b0111; // x=18, y=10
        pixel_data[10][19] = 4'b0111; // x=19, y=10
        pixel_data[10][20] = 4'b0111; // x=20, y=10
        pixel_data[10][21] = 4'b0111; // x=21, y=10
        pixel_data[10][22] = 4'b0111; // x=22, y=10
        pixel_data[10][23] = 4'b0111; // x=23, y=10
        pixel_data[10][24] = 4'b0111; // x=24, y=10
        pixel_data[10][25] = 4'b0111; // x=25, y=10
        pixel_data[10][26] = 4'b0111; // x=26, y=10
        pixel_data[10][27] = 4'b0111; // x=27, y=10
        pixel_data[10][28] = 4'b0111; // x=28, y=10
        pixel_data[10][29] = 4'b0111; // x=29, y=10
        pixel_data[10][30] = 4'b0111; // x=30, y=10
        pixel_data[10][31] = 4'b0111; // x=31, y=10
        pixel_data[10][32] = 4'b0111; // x=32, y=10
        pixel_data[10][33] = 4'b0111; // x=33, y=10
        pixel_data[10][34] = 4'b0111; // x=34, y=10
        pixel_data[10][35] = 4'b0111; // x=35, y=10
        pixel_data[10][36] = 4'b0111; // x=36, y=10
        pixel_data[10][37] = 4'b0111; // x=37, y=10
        pixel_data[10][38] = 4'b0111; // x=38, y=10
        pixel_data[10][39] = 4'b0111; // x=39, y=10
        pixel_data[10][40] = 4'b0111; // x=40, y=10
        pixel_data[10][41] = 4'b0111; // x=41, y=10
        pixel_data[10][42] = 4'b0111; // x=42, y=10
        pixel_data[10][43] = 4'b0111; // x=43, y=10
        pixel_data[10][44] = 4'b0111; // x=44, y=10
        pixel_data[10][45] = 4'b0111; // x=45, y=10
        pixel_data[10][46] = 4'b0111; // x=46, y=10
        pixel_data[10][47] = 4'b0111; // x=47, y=10
        pixel_data[10][48] = 4'b0111; // x=48, y=10
        pixel_data[10][49] = 4'b0111; // x=49, y=10
        pixel_data[10][50] = 4'b0111; // x=50, y=10
        pixel_data[10][51] = 4'b0111; // x=51, y=10
        pixel_data[10][52] = 4'b0111; // x=52, y=10
        pixel_data[10][53] = 4'b0111; // x=53, y=10
        pixel_data[10][54] = 4'b0111; // x=54, y=10
        pixel_data[10][55] = 4'b0111; // x=55, y=10
        pixel_data[10][56] = 4'b0111; // x=56, y=10
        pixel_data[10][57] = 4'b0111; // x=57, y=10
        pixel_data[10][58] = 4'b0111; // x=58, y=10
        pixel_data[10][59] = 4'b0111; // x=59, y=10
        pixel_data[10][60] = 4'b0111; // x=60, y=10
        pixel_data[10][61] = 4'b0111; // x=61, y=10
        pixel_data[10][62] = 4'b0111; // x=62, y=10
        pixel_data[10][63] = 4'b0111; // x=63, y=10
        pixel_data[10][64] = 4'b0111; // x=64, y=10
        pixel_data[10][65] = 4'b0111; // x=65, y=10
        pixel_data[10][66] = 4'b0111; // x=66, y=10
        pixel_data[10][67] = 4'b0111; // x=67, y=10
        pixel_data[10][68] = 4'b0111; // x=68, y=10
        pixel_data[10][69] = 4'b0111; // x=69, y=10
        pixel_data[10][70] = 4'b0111; // x=70, y=10
        pixel_data[10][71] = 4'b0111; // x=71, y=10
        pixel_data[10][72] = 4'b0111; // x=72, y=10
        pixel_data[10][73] = 4'b0111; // x=73, y=10
        pixel_data[10][74] = 4'b0111; // x=74, y=10
        pixel_data[10][75] = 4'b0111; // x=75, y=10
        pixel_data[10][76] = 4'b0111; // x=76, y=10
        pixel_data[10][77] = 4'b0111; // x=77, y=10
        pixel_data[10][78] = 4'b0111; // x=78, y=10
        pixel_data[10][79] = 4'b0111; // x=79, y=10
        pixel_data[10][80] = 4'b0111; // x=80, y=10
        pixel_data[10][81] = 4'b0111; // x=81, y=10
        pixel_data[10][82] = 4'b0111; // x=82, y=10
        pixel_data[10][83] = 4'b0111; // x=83, y=10
        pixel_data[10][84] = 4'b0111; // x=84, y=10
        pixel_data[10][85] = 4'b0111; // x=85, y=10
        pixel_data[10][86] = 4'b0111; // x=86, y=10
        pixel_data[10][87] = 4'b0111; // x=87, y=10
        pixel_data[10][88] = 4'b0111; // x=88, y=10
        pixel_data[10][89] = 4'b0111; // x=89, y=10
        pixel_data[10][90] = 4'b0111; // x=90, y=10
        pixel_data[10][91] = 4'b0111; // x=91, y=10
        pixel_data[10][92] = 4'b0111; // x=92, y=10
        pixel_data[10][93] = 4'b0111; // x=93, y=10
        pixel_data[10][94] = 4'b0111; // x=94, y=10
        pixel_data[10][95] = 4'b0111; // x=95, y=10
        pixel_data[10][96] = 4'b0111; // x=96, y=10
        pixel_data[10][97] = 4'b0111; // x=97, y=10
        pixel_data[10][98] = 4'b0111; // x=98, y=10
        pixel_data[10][99] = 4'b0111; // x=99, y=10
        pixel_data[10][100] = 4'b0111; // x=100, y=10
        pixel_data[10][101] = 4'b0111; // x=101, y=10
        pixel_data[10][102] = 4'b0111; // x=102, y=10
        pixel_data[10][103] = 4'b0111; // x=103, y=10
        pixel_data[10][104] = 4'b0111; // x=104, y=10
        pixel_data[10][105] = 4'b0111; // x=105, y=10
        pixel_data[10][106] = 4'b0111; // x=106, y=10
        pixel_data[10][107] = 4'b0111; // x=107, y=10
        pixel_data[10][108] = 4'b0111; // x=108, y=10
        pixel_data[10][109] = 4'b0111; // x=109, y=10
        pixel_data[10][110] = 4'b0111; // x=110, y=10
        pixel_data[10][111] = 4'b0111; // x=111, y=10
        pixel_data[10][112] = 4'b0111; // x=112, y=10
        pixel_data[10][113] = 4'b0111; // x=113, y=10
        pixel_data[10][114] = 4'b0111; // x=114, y=10
        pixel_data[10][115] = 4'b0111; // x=115, y=10
        pixel_data[10][116] = 4'b0111; // x=116, y=10
        pixel_data[10][117] = 4'b0111; // x=117, y=10
        pixel_data[10][118] = 4'b0111; // x=118, y=10
        pixel_data[10][119] = 4'b0111; // x=119, y=10
        pixel_data[10][120] = 4'b0111; // x=120, y=10
        pixel_data[10][121] = 4'b0111; // x=121, y=10
        pixel_data[10][122] = 4'b0111; // x=122, y=10
        pixel_data[10][123] = 4'b0111; // x=123, y=10
        pixel_data[10][124] = 4'b0111; // x=124, y=10
        pixel_data[10][125] = 4'b0111; // x=125, y=10
        pixel_data[10][126] = 4'b0111; // x=126, y=10
        pixel_data[10][127] = 4'b0111; // x=127, y=10
        pixel_data[10][128] = 4'b0111; // x=128, y=10
        pixel_data[10][129] = 4'b0111; // x=129, y=10
        pixel_data[10][130] = 4'b0111; // x=130, y=10
        pixel_data[10][131] = 4'b0111; // x=131, y=10
        pixel_data[10][132] = 4'b0111; // x=132, y=10
        pixel_data[10][133] = 4'b0111; // x=133, y=10
        pixel_data[10][134] = 4'b0111; // x=134, y=10
        pixel_data[10][135] = 4'b0111; // x=135, y=10
        pixel_data[10][136] = 4'b0111; // x=136, y=10
        pixel_data[10][137] = 4'b0111; // x=137, y=10
        pixel_data[10][138] = 4'b0111; // x=138, y=10
        pixel_data[10][139] = 4'b0111; // x=139, y=10
        pixel_data[10][140] = 4'b0111; // x=140, y=10
        pixel_data[10][141] = 4'b0111; // x=141, y=10
        pixel_data[10][142] = 4'b0111; // x=142, y=10
        pixel_data[10][143] = 4'b0111; // x=143, y=10
        pixel_data[10][144] = 4'b0111; // x=144, y=10
        pixel_data[10][145] = 4'b0111; // x=145, y=10
        pixel_data[10][146] = 4'b0111; // x=146, y=10
        pixel_data[10][147] = 4'b0111; // x=147, y=10
        pixel_data[10][148] = 4'b0111; // x=148, y=10
        pixel_data[10][149] = 4'b0111; // x=149, y=10
        pixel_data[10][150] = 4'b0111; // x=150, y=10
        pixel_data[10][151] = 4'b0111; // x=151, y=10
        pixel_data[10][152] = 4'b0111; // x=152, y=10
        pixel_data[10][153] = 4'b0111; // x=153, y=10
        pixel_data[10][154] = 4'b0111; // x=154, y=10
        pixel_data[10][155] = 4'b0111; // x=155, y=10
        pixel_data[10][156] = 4'b0111; // x=156, y=10
        pixel_data[10][157] = 4'b0111; // x=157, y=10
        pixel_data[10][158] = 4'b0111; // x=158, y=10
        pixel_data[10][159] = 4'b0111; // x=159, y=10
        pixel_data[10][160] = 4'b0111; // x=160, y=10
        pixel_data[10][161] = 4'b0111; // x=161, y=10
        pixel_data[10][162] = 4'b0111; // x=162, y=10
        pixel_data[10][163] = 4'b0111; // x=163, y=10
        pixel_data[10][164] = 4'b0111; // x=164, y=10
        pixel_data[10][165] = 4'b0111; // x=165, y=10
        pixel_data[10][166] = 4'b0111; // x=166, y=10
        pixel_data[10][167] = 4'b0111; // x=167, y=10
        pixel_data[10][168] = 4'b0111; // x=168, y=10
        pixel_data[10][169] = 4'b0111; // x=169, y=10
        pixel_data[10][170] = 4'b0111; // x=170, y=10
        pixel_data[10][171] = 4'b0111; // x=171, y=10
        pixel_data[10][172] = 4'b0111; // x=172, y=10
        pixel_data[10][173] = 4'b0111; // x=173, y=10
        pixel_data[10][174] = 4'b0111; // x=174, y=10
        pixel_data[10][175] = 4'b0111; // x=175, y=10
        pixel_data[10][176] = 4'b0111; // x=176, y=10
        pixel_data[10][177] = 4'b0111; // x=177, y=10
        pixel_data[10][178] = 4'b0111; // x=178, y=10
        pixel_data[10][179] = 4'b0111; // x=179, y=10
        pixel_data[11][0] = 4'b0111; // x=0, y=11
        pixel_data[11][1] = 4'b0111; // x=1, y=11
        pixel_data[11][2] = 4'b0111; // x=2, y=11
        pixel_data[11][3] = 4'b0111; // x=3, y=11
        pixel_data[11][4] = 4'b0111; // x=4, y=11
        pixel_data[11][5] = 4'b0111; // x=5, y=11
        pixel_data[11][6] = 4'b0111; // x=6, y=11
        pixel_data[11][7] = 4'b0111; // x=7, y=11
        pixel_data[11][8] = 4'b0111; // x=8, y=11
        pixel_data[11][9] = 4'b0111; // x=9, y=11
        pixel_data[11][10] = 4'b0111; // x=10, y=11
        pixel_data[11][11] = 4'b0111; // x=11, y=11
        pixel_data[11][12] = 4'b0111; // x=12, y=11
        pixel_data[11][13] = 4'b0111; // x=13, y=11
        pixel_data[11][14] = 4'b0111; // x=14, y=11
        pixel_data[11][15] = 4'b0111; // x=15, y=11
        pixel_data[11][16] = 4'b0111; // x=16, y=11
        pixel_data[11][17] = 4'b0111; // x=17, y=11
        pixel_data[11][18] = 4'b0111; // x=18, y=11
        pixel_data[11][19] = 4'b0111; // x=19, y=11
        pixel_data[11][20] = 4'b0111; // x=20, y=11
        pixel_data[11][21] = 4'b0111; // x=21, y=11
        pixel_data[11][22] = 4'b0111; // x=22, y=11
        pixel_data[11][23] = 4'b0111; // x=23, y=11
        pixel_data[11][24] = 4'b0111; // x=24, y=11
        pixel_data[11][25] = 4'b0111; // x=25, y=11
        pixel_data[11][26] = 4'b0111; // x=26, y=11
        pixel_data[11][27] = 4'b0111; // x=27, y=11
        pixel_data[11][28] = 4'b0111; // x=28, y=11
        pixel_data[11][29] = 4'b0111; // x=29, y=11
        pixel_data[11][30] = 4'b0111; // x=30, y=11
        pixel_data[11][31] = 4'b0111; // x=31, y=11
        pixel_data[11][32] = 4'b0111; // x=32, y=11
        pixel_data[11][33] = 4'b0111; // x=33, y=11
        pixel_data[11][34] = 4'b0111; // x=34, y=11
        pixel_data[11][35] = 4'b0111; // x=35, y=11
        pixel_data[11][36] = 4'b0111; // x=36, y=11
        pixel_data[11][37] = 4'b0111; // x=37, y=11
        pixel_data[11][38] = 4'b0111; // x=38, y=11
        pixel_data[11][39] = 4'b0111; // x=39, y=11
        pixel_data[11][40] = 4'b0111; // x=40, y=11
        pixel_data[11][41] = 4'b0111; // x=41, y=11
        pixel_data[11][42] = 4'b0111; // x=42, y=11
        pixel_data[11][43] = 4'b0111; // x=43, y=11
        pixel_data[11][44] = 4'b0111; // x=44, y=11
        pixel_data[11][45] = 4'b0111; // x=45, y=11
        pixel_data[11][46] = 4'b0111; // x=46, y=11
        pixel_data[11][47] = 4'b0111; // x=47, y=11
        pixel_data[11][48] = 4'b0111; // x=48, y=11
        pixel_data[11][49] = 4'b0111; // x=49, y=11
        pixel_data[11][50] = 4'b0111; // x=50, y=11
        pixel_data[11][51] = 4'b0111; // x=51, y=11
        pixel_data[11][52] = 4'b0111; // x=52, y=11
        pixel_data[11][53] = 4'b0111; // x=53, y=11
        pixel_data[11][54] = 4'b0111; // x=54, y=11
        pixel_data[11][55] = 4'b0111; // x=55, y=11
        pixel_data[11][56] = 4'b0111; // x=56, y=11
        pixel_data[11][57] = 4'b0111; // x=57, y=11
        pixel_data[11][58] = 4'b0111; // x=58, y=11
        pixel_data[11][59] = 4'b0111; // x=59, y=11
        pixel_data[11][60] = 4'b0111; // x=60, y=11
        pixel_data[11][61] = 4'b0111; // x=61, y=11
        pixel_data[11][62] = 4'b0111; // x=62, y=11
        pixel_data[11][63] = 4'b0111; // x=63, y=11
        pixel_data[11][64] = 4'b0111; // x=64, y=11
        pixel_data[11][65] = 4'b0111; // x=65, y=11
        pixel_data[11][66] = 4'b0111; // x=66, y=11
        pixel_data[11][67] = 4'b0111; // x=67, y=11
        pixel_data[11][68] = 4'b0111; // x=68, y=11
        pixel_data[11][69] = 4'b0111; // x=69, y=11
        pixel_data[11][70] = 4'b0111; // x=70, y=11
        pixel_data[11][71] = 4'b0111; // x=71, y=11
        pixel_data[11][72] = 4'b0111; // x=72, y=11
        pixel_data[11][73] = 4'b0111; // x=73, y=11
        pixel_data[11][74] = 4'b0111; // x=74, y=11
        pixel_data[11][75] = 4'b0111; // x=75, y=11
        pixel_data[11][76] = 4'b0111; // x=76, y=11
        pixel_data[11][77] = 4'b0111; // x=77, y=11
        pixel_data[11][78] = 4'b0111; // x=78, y=11
        pixel_data[11][79] = 4'b0111; // x=79, y=11
        pixel_data[11][80] = 4'b0111; // x=80, y=11
        pixel_data[11][81] = 4'b0111; // x=81, y=11
        pixel_data[11][82] = 4'b0111; // x=82, y=11
        pixel_data[11][83] = 4'b0111; // x=83, y=11
        pixel_data[11][84] = 4'b0111; // x=84, y=11
        pixel_data[11][85] = 4'b0111; // x=85, y=11
        pixel_data[11][86] = 4'b0111; // x=86, y=11
        pixel_data[11][87] = 4'b0111; // x=87, y=11
        pixel_data[11][88] = 4'b0111; // x=88, y=11
        pixel_data[11][89] = 4'b0111; // x=89, y=11
        pixel_data[11][90] = 4'b0111; // x=90, y=11
        pixel_data[11][91] = 4'b0111; // x=91, y=11
        pixel_data[11][92] = 4'b0111; // x=92, y=11
        pixel_data[11][93] = 4'b0111; // x=93, y=11
        pixel_data[11][94] = 4'b0111; // x=94, y=11
        pixel_data[11][95] = 4'b0111; // x=95, y=11
        pixel_data[11][96] = 4'b0111; // x=96, y=11
        pixel_data[11][97] = 4'b0111; // x=97, y=11
        pixel_data[11][98] = 4'b0111; // x=98, y=11
        pixel_data[11][99] = 4'b0111; // x=99, y=11
        pixel_data[11][100] = 4'b0111; // x=100, y=11
        pixel_data[11][101] = 4'b0111; // x=101, y=11
        pixel_data[11][102] = 4'b0111; // x=102, y=11
        pixel_data[11][103] = 4'b0111; // x=103, y=11
        pixel_data[11][104] = 4'b0111; // x=104, y=11
        pixel_data[11][105] = 4'b0111; // x=105, y=11
        pixel_data[11][106] = 4'b0111; // x=106, y=11
        pixel_data[11][107] = 4'b0111; // x=107, y=11
        pixel_data[11][108] = 4'b0111; // x=108, y=11
        pixel_data[11][109] = 4'b0111; // x=109, y=11
        pixel_data[11][110] = 4'b0111; // x=110, y=11
        pixel_data[11][111] = 4'b0111; // x=111, y=11
        pixel_data[11][112] = 4'b0111; // x=112, y=11
        pixel_data[11][113] = 4'b0111; // x=113, y=11
        pixel_data[11][114] = 4'b0111; // x=114, y=11
        pixel_data[11][115] = 4'b0111; // x=115, y=11
        pixel_data[11][116] = 4'b0111; // x=116, y=11
        pixel_data[11][117] = 4'b0111; // x=117, y=11
        pixel_data[11][118] = 4'b0111; // x=118, y=11
        pixel_data[11][119] = 4'b0111; // x=119, y=11
        pixel_data[11][120] = 4'b0111; // x=120, y=11
        pixel_data[11][121] = 4'b0111; // x=121, y=11
        pixel_data[11][122] = 4'b0111; // x=122, y=11
        pixel_data[11][123] = 4'b0111; // x=123, y=11
        pixel_data[11][124] = 4'b0111; // x=124, y=11
        pixel_data[11][125] = 4'b0111; // x=125, y=11
        pixel_data[11][126] = 4'b0111; // x=126, y=11
        pixel_data[11][127] = 4'b0111; // x=127, y=11
        pixel_data[11][128] = 4'b0111; // x=128, y=11
        pixel_data[11][129] = 4'b0111; // x=129, y=11
        pixel_data[11][130] = 4'b0111; // x=130, y=11
        pixel_data[11][131] = 4'b0111; // x=131, y=11
        pixel_data[11][132] = 4'b0111; // x=132, y=11
        pixel_data[11][133] = 4'b0111; // x=133, y=11
        pixel_data[11][134] = 4'b0111; // x=134, y=11
        pixel_data[11][135] = 4'b0111; // x=135, y=11
        pixel_data[11][136] = 4'b0111; // x=136, y=11
        pixel_data[11][137] = 4'b0111; // x=137, y=11
        pixel_data[11][138] = 4'b0111; // x=138, y=11
        pixel_data[11][139] = 4'b0111; // x=139, y=11
        pixel_data[11][140] = 4'b0111; // x=140, y=11
        pixel_data[11][141] = 4'b0111; // x=141, y=11
        pixel_data[11][142] = 4'b0111; // x=142, y=11
        pixel_data[11][143] = 4'b0111; // x=143, y=11
        pixel_data[11][144] = 4'b0111; // x=144, y=11
        pixel_data[11][145] = 4'b0111; // x=145, y=11
        pixel_data[11][146] = 4'b0111; // x=146, y=11
        pixel_data[11][147] = 4'b0111; // x=147, y=11
        pixel_data[11][148] = 4'b0111; // x=148, y=11
        pixel_data[11][149] = 4'b0111; // x=149, y=11
        pixel_data[11][150] = 4'b0111; // x=150, y=11
        pixel_data[11][151] = 4'b0111; // x=151, y=11
        pixel_data[11][152] = 4'b0111; // x=152, y=11
        pixel_data[11][153] = 4'b0111; // x=153, y=11
        pixel_data[11][154] = 4'b0111; // x=154, y=11
        pixel_data[11][155] = 4'b0111; // x=155, y=11
        pixel_data[11][156] = 4'b0111; // x=156, y=11
        pixel_data[11][157] = 4'b0111; // x=157, y=11
        pixel_data[11][158] = 4'b0111; // x=158, y=11
        pixel_data[11][159] = 4'b0111; // x=159, y=11
        pixel_data[11][160] = 4'b0111; // x=160, y=11
        pixel_data[11][161] = 4'b0111; // x=161, y=11
        pixel_data[11][162] = 4'b0111; // x=162, y=11
        pixel_data[11][163] = 4'b0111; // x=163, y=11
        pixel_data[11][164] = 4'b0111; // x=164, y=11
        pixel_data[11][165] = 4'b0111; // x=165, y=11
        pixel_data[11][166] = 4'b0111; // x=166, y=11
        pixel_data[11][167] = 4'b0111; // x=167, y=11
        pixel_data[11][168] = 4'b0111; // x=168, y=11
        pixel_data[11][169] = 4'b0111; // x=169, y=11
        pixel_data[11][170] = 4'b0111; // x=170, y=11
        pixel_data[11][171] = 4'b0111; // x=171, y=11
        pixel_data[11][172] = 4'b0111; // x=172, y=11
        pixel_data[11][173] = 4'b0111; // x=173, y=11
        pixel_data[11][174] = 4'b0111; // x=174, y=11
        pixel_data[11][175] = 4'b0111; // x=175, y=11
        pixel_data[11][176] = 4'b0111; // x=176, y=11
        pixel_data[11][177] = 4'b0111; // x=177, y=11
        pixel_data[11][178] = 4'b0111; // x=178, y=11
        pixel_data[11][179] = 4'b0111; // x=179, y=11
        pixel_data[12][0] = 4'b0111; // x=0, y=12
        pixel_data[12][1] = 4'b0111; // x=1, y=12
        pixel_data[12][2] = 4'b0111; // x=2, y=12
        pixel_data[12][3] = 4'b0111; // x=3, y=12
        pixel_data[12][4] = 4'b0111; // x=4, y=12
        pixel_data[12][5] = 4'b0111; // x=5, y=12
        pixel_data[12][6] = 4'b0111; // x=6, y=12
        pixel_data[12][7] = 4'b0111; // x=7, y=12
        pixel_data[12][8] = 4'b0111; // x=8, y=12
        pixel_data[12][9] = 4'b0111; // x=9, y=12
        pixel_data[12][10] = 4'b0111; // x=10, y=12
        pixel_data[12][11] = 4'b0111; // x=11, y=12
        pixel_data[12][12] = 4'b0111; // x=12, y=12
        pixel_data[12][13] = 4'b0111; // x=13, y=12
        pixel_data[12][14] = 4'b0111; // x=14, y=12
        pixel_data[12][15] = 4'b0111; // x=15, y=12
        pixel_data[12][16] = 4'b0111; // x=16, y=12
        pixel_data[12][17] = 4'b0111; // x=17, y=12
        pixel_data[12][18] = 4'b0111; // x=18, y=12
        pixel_data[12][19] = 4'b0111; // x=19, y=12
        pixel_data[12][20] = 4'b0111; // x=20, y=12
        pixel_data[12][21] = 4'b0111; // x=21, y=12
        pixel_data[12][22] = 4'b0111; // x=22, y=12
        pixel_data[12][23] = 4'b0111; // x=23, y=12
        pixel_data[12][24] = 4'b0111; // x=24, y=12
        pixel_data[12][25] = 4'b0111; // x=25, y=12
        pixel_data[12][26] = 4'b0111; // x=26, y=12
        pixel_data[12][27] = 4'b0111; // x=27, y=12
        pixel_data[12][28] = 4'b0111; // x=28, y=12
        pixel_data[12][29] = 4'b0111; // x=29, y=12
        pixel_data[12][30] = 4'b0111; // x=30, y=12
        pixel_data[12][31] = 4'b0111; // x=31, y=12
        pixel_data[12][32] = 4'b0111; // x=32, y=12
        pixel_data[12][33] = 4'b0111; // x=33, y=12
        pixel_data[12][34] = 4'b0111; // x=34, y=12
        pixel_data[12][35] = 4'b0111; // x=35, y=12
        pixel_data[12][36] = 4'b0111; // x=36, y=12
        pixel_data[12][37] = 4'b0111; // x=37, y=12
        pixel_data[12][38] = 4'b0111; // x=38, y=12
        pixel_data[12][39] = 4'b0111; // x=39, y=12
        pixel_data[12][40] = 4'b0111; // x=40, y=12
        pixel_data[12][41] = 4'b0111; // x=41, y=12
        pixel_data[12][42] = 4'b0111; // x=42, y=12
        pixel_data[12][43] = 4'b0111; // x=43, y=12
        pixel_data[12][44] = 4'b0111; // x=44, y=12
        pixel_data[12][45] = 4'b0111; // x=45, y=12
        pixel_data[12][46] = 4'b0111; // x=46, y=12
        pixel_data[12][47] = 4'b0111; // x=47, y=12
        pixel_data[12][48] = 4'b0111; // x=48, y=12
        pixel_data[12][49] = 4'b0111; // x=49, y=12
        pixel_data[12][50] = 4'b0111; // x=50, y=12
        pixel_data[12][51] = 4'b0111; // x=51, y=12
        pixel_data[12][52] = 4'b0111; // x=52, y=12
        pixel_data[12][53] = 4'b0111; // x=53, y=12
        pixel_data[12][54] = 4'b0111; // x=54, y=12
        pixel_data[12][55] = 4'b0111; // x=55, y=12
        pixel_data[12][56] = 4'b0111; // x=56, y=12
        pixel_data[12][57] = 4'b0111; // x=57, y=12
        pixel_data[12][58] = 4'b0111; // x=58, y=12
        pixel_data[12][59] = 4'b0111; // x=59, y=12
        pixel_data[12][60] = 4'b0111; // x=60, y=12
        pixel_data[12][61] = 4'b0111; // x=61, y=12
        pixel_data[12][62] = 4'b0111; // x=62, y=12
        pixel_data[12][63] = 4'b0111; // x=63, y=12
        pixel_data[12][64] = 4'b0111; // x=64, y=12
        pixel_data[12][65] = 4'b0111; // x=65, y=12
        pixel_data[12][66] = 4'b0111; // x=66, y=12
        pixel_data[12][67] = 4'b0111; // x=67, y=12
        pixel_data[12][68] = 4'b0111; // x=68, y=12
        pixel_data[12][69] = 4'b0111; // x=69, y=12
        pixel_data[12][70] = 4'b0111; // x=70, y=12
        pixel_data[12][71] = 4'b0111; // x=71, y=12
        pixel_data[12][72] = 4'b0111; // x=72, y=12
        pixel_data[12][73] = 4'b0111; // x=73, y=12
        pixel_data[12][74] = 4'b0111; // x=74, y=12
        pixel_data[12][75] = 4'b0111; // x=75, y=12
        pixel_data[12][76] = 4'b0111; // x=76, y=12
        pixel_data[12][77] = 4'b0111; // x=77, y=12
        pixel_data[12][78] = 4'b0111; // x=78, y=12
        pixel_data[12][79] = 4'b0111; // x=79, y=12
        pixel_data[12][80] = 4'b0111; // x=80, y=12
        pixel_data[12][81] = 4'b0111; // x=81, y=12
        pixel_data[12][82] = 4'b0111; // x=82, y=12
        pixel_data[12][83] = 4'b0111; // x=83, y=12
        pixel_data[12][84] = 4'b0111; // x=84, y=12
        pixel_data[12][85] = 4'b0111; // x=85, y=12
        pixel_data[12][86] = 4'b0111; // x=86, y=12
        pixel_data[12][87] = 4'b0111; // x=87, y=12
        pixel_data[12][88] = 4'b0111; // x=88, y=12
        pixel_data[12][89] = 4'b0111; // x=89, y=12
        pixel_data[12][90] = 4'b0111; // x=90, y=12
        pixel_data[12][91] = 4'b0111; // x=91, y=12
        pixel_data[12][92] = 4'b0111; // x=92, y=12
        pixel_data[12][93] = 4'b0111; // x=93, y=12
        pixel_data[12][94] = 4'b0111; // x=94, y=12
        pixel_data[12][95] = 4'b0111; // x=95, y=12
        pixel_data[12][96] = 4'b0111; // x=96, y=12
        pixel_data[12][97] = 4'b0111; // x=97, y=12
        pixel_data[12][98] = 4'b0111; // x=98, y=12
        pixel_data[12][99] = 4'b0111; // x=99, y=12
        pixel_data[12][100] = 4'b0111; // x=100, y=12
        pixel_data[12][101] = 4'b0111; // x=101, y=12
        pixel_data[12][102] = 4'b0111; // x=102, y=12
        pixel_data[12][103] = 4'b0111; // x=103, y=12
        pixel_data[12][104] = 4'b0111; // x=104, y=12
        pixel_data[12][105] = 4'b0111; // x=105, y=12
        pixel_data[12][106] = 4'b0111; // x=106, y=12
        pixel_data[12][107] = 4'b0111; // x=107, y=12
        pixel_data[12][108] = 4'b0111; // x=108, y=12
        pixel_data[12][109] = 4'b0111; // x=109, y=12
        pixel_data[12][110] = 4'b0111; // x=110, y=12
        pixel_data[12][111] = 4'b0111; // x=111, y=12
        pixel_data[12][112] = 4'b0111; // x=112, y=12
        pixel_data[12][113] = 4'b0111; // x=113, y=12
        pixel_data[12][114] = 4'b0111; // x=114, y=12
        pixel_data[12][115] = 4'b0111; // x=115, y=12
        pixel_data[12][116] = 4'b0111; // x=116, y=12
        pixel_data[12][117] = 4'b0111; // x=117, y=12
        pixel_data[12][118] = 4'b0111; // x=118, y=12
        pixel_data[12][119] = 4'b0111; // x=119, y=12
        pixel_data[12][120] = 4'b0111; // x=120, y=12
        pixel_data[12][121] = 4'b0111; // x=121, y=12
        pixel_data[12][122] = 4'b0111; // x=122, y=12
        pixel_data[12][123] = 4'b0111; // x=123, y=12
        pixel_data[12][124] = 4'b0111; // x=124, y=12
        pixel_data[12][125] = 4'b0111; // x=125, y=12
        pixel_data[12][126] = 4'b0111; // x=126, y=12
        pixel_data[12][127] = 4'b0111; // x=127, y=12
        pixel_data[12][128] = 4'b0111; // x=128, y=12
        pixel_data[12][129] = 4'b0111; // x=129, y=12
        pixel_data[12][130] = 4'b0111; // x=130, y=12
        pixel_data[12][131] = 4'b0111; // x=131, y=12
        pixel_data[12][132] = 4'b0111; // x=132, y=12
        pixel_data[12][133] = 4'b0111; // x=133, y=12
        pixel_data[12][134] = 4'b0111; // x=134, y=12
        pixel_data[12][135] = 4'b0111; // x=135, y=12
        pixel_data[12][136] = 4'b0111; // x=136, y=12
        pixel_data[12][137] = 4'b0111; // x=137, y=12
        pixel_data[12][138] = 4'b0111; // x=138, y=12
        pixel_data[12][139] = 4'b0111; // x=139, y=12
        pixel_data[12][140] = 4'b0111; // x=140, y=12
        pixel_data[12][141] = 4'b0111; // x=141, y=12
        pixel_data[12][142] = 4'b0111; // x=142, y=12
        pixel_data[12][143] = 4'b0111; // x=143, y=12
        pixel_data[12][144] = 4'b0111; // x=144, y=12
        pixel_data[12][145] = 4'b0111; // x=145, y=12
        pixel_data[12][146] = 4'b0111; // x=146, y=12
        pixel_data[12][147] = 4'b0111; // x=147, y=12
        pixel_data[12][148] = 4'b0111; // x=148, y=12
        pixel_data[12][149] = 4'b0111; // x=149, y=12
        pixel_data[12][150] = 4'b0111; // x=150, y=12
        pixel_data[12][151] = 4'b0111; // x=151, y=12
        pixel_data[12][152] = 4'b0111; // x=152, y=12
        pixel_data[12][153] = 4'b0111; // x=153, y=12
        pixel_data[12][154] = 4'b0111; // x=154, y=12
        pixel_data[12][155] = 4'b0111; // x=155, y=12
        pixel_data[12][156] = 4'b0111; // x=156, y=12
        pixel_data[12][157] = 4'b0111; // x=157, y=12
        pixel_data[12][158] = 4'b0111; // x=158, y=12
        pixel_data[12][159] = 4'b0111; // x=159, y=12
        pixel_data[12][160] = 4'b0111; // x=160, y=12
        pixel_data[12][161] = 4'b0111; // x=161, y=12
        pixel_data[12][162] = 4'b0111; // x=162, y=12
        pixel_data[12][163] = 4'b0111; // x=163, y=12
        pixel_data[12][164] = 4'b0111; // x=164, y=12
        pixel_data[12][165] = 4'b0111; // x=165, y=12
        pixel_data[12][166] = 4'b0111; // x=166, y=12
        pixel_data[12][167] = 4'b0111; // x=167, y=12
        pixel_data[12][168] = 4'b0111; // x=168, y=12
        pixel_data[12][169] = 4'b0111; // x=169, y=12
        pixel_data[12][170] = 4'b0111; // x=170, y=12
        pixel_data[12][171] = 4'b0111; // x=171, y=12
        pixel_data[12][172] = 4'b0111; // x=172, y=12
        pixel_data[12][173] = 4'b0111; // x=173, y=12
        pixel_data[12][174] = 4'b0111; // x=174, y=12
        pixel_data[12][175] = 4'b0111; // x=175, y=12
        pixel_data[12][176] = 4'b0111; // x=176, y=12
        pixel_data[12][177] = 4'b0111; // x=177, y=12
        pixel_data[12][178] = 4'b0111; // x=178, y=12
        pixel_data[12][179] = 4'b0111; // x=179, y=12
        pixel_data[13][0] = 4'b0111; // x=0, y=13
        pixel_data[13][1] = 4'b0111; // x=1, y=13
        pixel_data[13][2] = 4'b0111; // x=2, y=13
        pixel_data[13][3] = 4'b0111; // x=3, y=13
        pixel_data[13][4] = 4'b0111; // x=4, y=13
        pixel_data[13][5] = 4'b0111; // x=5, y=13
        pixel_data[13][6] = 4'b0111; // x=6, y=13
        pixel_data[13][7] = 4'b0111; // x=7, y=13
        pixel_data[13][8] = 4'b0111; // x=8, y=13
        pixel_data[13][9] = 4'b0111; // x=9, y=13
        pixel_data[13][10] = 4'b0111; // x=10, y=13
        pixel_data[13][11] = 4'b0111; // x=11, y=13
        pixel_data[13][12] = 4'b0111; // x=12, y=13
        pixel_data[13][13] = 4'b0111; // x=13, y=13
        pixel_data[13][14] = 4'b0111; // x=14, y=13
        pixel_data[13][15] = 4'b0111; // x=15, y=13
        pixel_data[13][16] = 4'b0111; // x=16, y=13
        pixel_data[13][17] = 4'b0111; // x=17, y=13
        pixel_data[13][18] = 4'b0111; // x=18, y=13
        pixel_data[13][19] = 4'b0111; // x=19, y=13
        pixel_data[13][20] = 4'b0111; // x=20, y=13
        pixel_data[13][21] = 4'b0111; // x=21, y=13
        pixel_data[13][22] = 4'b0111; // x=22, y=13
        pixel_data[13][23] = 4'b0111; // x=23, y=13
        pixel_data[13][24] = 4'b0111; // x=24, y=13
        pixel_data[13][25] = 4'b0111; // x=25, y=13
        pixel_data[13][26] = 4'b0111; // x=26, y=13
        pixel_data[13][27] = 4'b0111; // x=27, y=13
        pixel_data[13][28] = 4'b0111; // x=28, y=13
        pixel_data[13][29] = 4'b0111; // x=29, y=13
        pixel_data[13][30] = 4'b0111; // x=30, y=13
        pixel_data[13][31] = 4'b0111; // x=31, y=13
        pixel_data[13][32] = 4'b0111; // x=32, y=13
        pixel_data[13][33] = 4'b0111; // x=33, y=13
        pixel_data[13][34] = 4'b0111; // x=34, y=13
        pixel_data[13][35] = 4'b0111; // x=35, y=13
        pixel_data[13][36] = 4'b0111; // x=36, y=13
        pixel_data[13][37] = 4'b0111; // x=37, y=13
        pixel_data[13][38] = 4'b0111; // x=38, y=13
        pixel_data[13][39] = 4'b0111; // x=39, y=13
        pixel_data[13][40] = 4'b0111; // x=40, y=13
        pixel_data[13][41] = 4'b0111; // x=41, y=13
        pixel_data[13][42] = 4'b0111; // x=42, y=13
        pixel_data[13][43] = 4'b0111; // x=43, y=13
        pixel_data[13][44] = 4'b0111; // x=44, y=13
        pixel_data[13][45] = 4'b0111; // x=45, y=13
        pixel_data[13][46] = 4'b0111; // x=46, y=13
        pixel_data[13][47] = 4'b0111; // x=47, y=13
        pixel_data[13][48] = 4'b0111; // x=48, y=13
        pixel_data[13][49] = 4'b0111; // x=49, y=13
        pixel_data[13][50] = 4'b0111; // x=50, y=13
        pixel_data[13][51] = 4'b0111; // x=51, y=13
        pixel_data[13][52] = 4'b0111; // x=52, y=13
        pixel_data[13][53] = 4'b0111; // x=53, y=13
        pixel_data[13][54] = 4'b0111; // x=54, y=13
        pixel_data[13][55] = 4'b0111; // x=55, y=13
        pixel_data[13][56] = 4'b0111; // x=56, y=13
        pixel_data[13][57] = 4'b0111; // x=57, y=13
        pixel_data[13][58] = 4'b0111; // x=58, y=13
        pixel_data[13][59] = 4'b0111; // x=59, y=13
        pixel_data[13][60] = 4'b0111; // x=60, y=13
        pixel_data[13][61] = 4'b0111; // x=61, y=13
        pixel_data[13][62] = 4'b0111; // x=62, y=13
        pixel_data[13][63] = 4'b0111; // x=63, y=13
        pixel_data[13][64] = 4'b0111; // x=64, y=13
        pixel_data[13][65] = 4'b0111; // x=65, y=13
        pixel_data[13][66] = 4'b0111; // x=66, y=13
        pixel_data[13][67] = 4'b0111; // x=67, y=13
        pixel_data[13][68] = 4'b0111; // x=68, y=13
        pixel_data[13][69] = 4'b0111; // x=69, y=13
        pixel_data[13][70] = 4'b0111; // x=70, y=13
        pixel_data[13][71] = 4'b0111; // x=71, y=13
        pixel_data[13][72] = 4'b0111; // x=72, y=13
        pixel_data[13][73] = 4'b0111; // x=73, y=13
        pixel_data[13][74] = 4'b0111; // x=74, y=13
        pixel_data[13][75] = 4'b0111; // x=75, y=13
        pixel_data[13][76] = 4'b0111; // x=76, y=13
        pixel_data[13][77] = 4'b0111; // x=77, y=13
        pixel_data[13][78] = 4'b0111; // x=78, y=13
        pixel_data[13][79] = 4'b0111; // x=79, y=13
        pixel_data[13][80] = 4'b0111; // x=80, y=13
        pixel_data[13][81] = 4'b0111; // x=81, y=13
        pixel_data[13][82] = 4'b0111; // x=82, y=13
        pixel_data[13][83] = 4'b0111; // x=83, y=13
        pixel_data[13][84] = 4'b0111; // x=84, y=13
        pixel_data[13][85] = 4'b0111; // x=85, y=13
        pixel_data[13][86] = 4'b0111; // x=86, y=13
        pixel_data[13][87] = 4'b0111; // x=87, y=13
        pixel_data[13][88] = 4'b0111; // x=88, y=13
        pixel_data[13][89] = 4'b0111; // x=89, y=13
        pixel_data[13][90] = 4'b0111; // x=90, y=13
        pixel_data[13][91] = 4'b0111; // x=91, y=13
        pixel_data[13][92] = 4'b0111; // x=92, y=13
        pixel_data[13][93] = 4'b0111; // x=93, y=13
        pixel_data[13][94] = 4'b0111; // x=94, y=13
        pixel_data[13][95] = 4'b0111; // x=95, y=13
        pixel_data[13][96] = 4'b0111; // x=96, y=13
        pixel_data[13][97] = 4'b0111; // x=97, y=13
        pixel_data[13][98] = 4'b0111; // x=98, y=13
        pixel_data[13][99] = 4'b0111; // x=99, y=13
        pixel_data[13][100] = 4'b0111; // x=100, y=13
        pixel_data[13][101] = 4'b0111; // x=101, y=13
        pixel_data[13][102] = 4'b0111; // x=102, y=13
        pixel_data[13][103] = 4'b0111; // x=103, y=13
        pixel_data[13][104] = 4'b0111; // x=104, y=13
        pixel_data[13][105] = 4'b0111; // x=105, y=13
        pixel_data[13][106] = 4'b0111; // x=106, y=13
        pixel_data[13][107] = 4'b0111; // x=107, y=13
        pixel_data[13][108] = 4'b0111; // x=108, y=13
        pixel_data[13][109] = 4'b0111; // x=109, y=13
        pixel_data[13][110] = 4'b0111; // x=110, y=13
        pixel_data[13][111] = 4'b0111; // x=111, y=13
        pixel_data[13][112] = 4'b0111; // x=112, y=13
        pixel_data[13][113] = 4'b0111; // x=113, y=13
        pixel_data[13][114] = 4'b0111; // x=114, y=13
        pixel_data[13][115] = 4'b0111; // x=115, y=13
        pixel_data[13][116] = 4'b0111; // x=116, y=13
        pixel_data[13][117] = 4'b0111; // x=117, y=13
        pixel_data[13][118] = 4'b0111; // x=118, y=13
        pixel_data[13][119] = 4'b0111; // x=119, y=13
        pixel_data[13][120] = 4'b0111; // x=120, y=13
        pixel_data[13][121] = 4'b0111; // x=121, y=13
        pixel_data[13][122] = 4'b0111; // x=122, y=13
        pixel_data[13][123] = 4'b0111; // x=123, y=13
        pixel_data[13][124] = 4'b0111; // x=124, y=13
        pixel_data[13][125] = 4'b0111; // x=125, y=13
        pixel_data[13][126] = 4'b0111; // x=126, y=13
        pixel_data[13][127] = 4'b0111; // x=127, y=13
        pixel_data[13][128] = 4'b0111; // x=128, y=13
        pixel_data[13][129] = 4'b0111; // x=129, y=13
        pixel_data[13][130] = 4'b0111; // x=130, y=13
        pixel_data[13][131] = 4'b0111; // x=131, y=13
        pixel_data[13][132] = 4'b0111; // x=132, y=13
        pixel_data[13][133] = 4'b0111; // x=133, y=13
        pixel_data[13][134] = 4'b0111; // x=134, y=13
        pixel_data[13][135] = 4'b0111; // x=135, y=13
        pixel_data[13][136] = 4'b0111; // x=136, y=13
        pixel_data[13][137] = 4'b0111; // x=137, y=13
        pixel_data[13][138] = 4'b0111; // x=138, y=13
        pixel_data[13][139] = 4'b0111; // x=139, y=13
        pixel_data[13][140] = 4'b0111; // x=140, y=13
        pixel_data[13][141] = 4'b0111; // x=141, y=13
        pixel_data[13][142] = 4'b0111; // x=142, y=13
        pixel_data[13][143] = 4'b0111; // x=143, y=13
        pixel_data[13][144] = 4'b0111; // x=144, y=13
        pixel_data[13][145] = 4'b0111; // x=145, y=13
        pixel_data[13][146] = 4'b0111; // x=146, y=13
        pixel_data[13][147] = 4'b0111; // x=147, y=13
        pixel_data[13][148] = 4'b0111; // x=148, y=13
        pixel_data[13][149] = 4'b0111; // x=149, y=13
        pixel_data[13][150] = 4'b0111; // x=150, y=13
        pixel_data[13][151] = 4'b0111; // x=151, y=13
        pixel_data[13][152] = 4'b0111; // x=152, y=13
        pixel_data[13][153] = 4'b0111; // x=153, y=13
        pixel_data[13][154] = 4'b0111; // x=154, y=13
        pixel_data[13][155] = 4'b0111; // x=155, y=13
        pixel_data[13][156] = 4'b0111; // x=156, y=13
        pixel_data[13][157] = 4'b0111; // x=157, y=13
        pixel_data[13][158] = 4'b0111; // x=158, y=13
        pixel_data[13][159] = 4'b0111; // x=159, y=13
        pixel_data[13][160] = 4'b0111; // x=160, y=13
        pixel_data[13][161] = 4'b0111; // x=161, y=13
        pixel_data[13][162] = 4'b0111; // x=162, y=13
        pixel_data[13][163] = 4'b0111; // x=163, y=13
        pixel_data[13][164] = 4'b0111; // x=164, y=13
        pixel_data[13][165] = 4'b0111; // x=165, y=13
        pixel_data[13][166] = 4'b0111; // x=166, y=13
        pixel_data[13][167] = 4'b0111; // x=167, y=13
        pixel_data[13][168] = 4'b0111; // x=168, y=13
        pixel_data[13][169] = 4'b0111; // x=169, y=13
        pixel_data[13][170] = 4'b0111; // x=170, y=13
        pixel_data[13][171] = 4'b0111; // x=171, y=13
        pixel_data[13][172] = 4'b0111; // x=172, y=13
        pixel_data[13][173] = 4'b0111; // x=173, y=13
        pixel_data[13][174] = 4'b0111; // x=174, y=13
        pixel_data[13][175] = 4'b0111; // x=175, y=13
        pixel_data[13][176] = 4'b0111; // x=176, y=13
        pixel_data[13][177] = 4'b0111; // x=177, y=13
        pixel_data[13][178] = 4'b0111; // x=178, y=13
        pixel_data[13][179] = 4'b0111; // x=179, y=13
        pixel_data[14][0] = 4'b0111; // x=0, y=14
        pixel_data[14][1] = 4'b0111; // x=1, y=14
        pixel_data[14][2] = 4'b0111; // x=2, y=14
        pixel_data[14][3] = 4'b0111; // x=3, y=14
        pixel_data[14][4] = 4'b0111; // x=4, y=14
        pixel_data[14][5] = 4'b0111; // x=5, y=14
        pixel_data[14][6] = 4'b0111; // x=6, y=14
        pixel_data[14][7] = 4'b0111; // x=7, y=14
        pixel_data[14][8] = 4'b0111; // x=8, y=14
        pixel_data[14][9] = 4'b0111; // x=9, y=14
        pixel_data[14][10] = 4'b0111; // x=10, y=14
        pixel_data[14][11] = 4'b0111; // x=11, y=14
        pixel_data[14][12] = 4'b0111; // x=12, y=14
        pixel_data[14][13] = 4'b0111; // x=13, y=14
        pixel_data[14][14] = 4'b0111; // x=14, y=14
        pixel_data[14][15] = 4'b0111; // x=15, y=14
        pixel_data[14][16] = 4'b0111; // x=16, y=14
        pixel_data[14][17] = 4'b0111; // x=17, y=14
        pixel_data[14][18] = 4'b0111; // x=18, y=14
        pixel_data[14][19] = 4'b0111; // x=19, y=14
        pixel_data[14][20] = 4'b0111; // x=20, y=14
        pixel_data[14][21] = 4'b0111; // x=21, y=14
        pixel_data[14][22] = 4'b0000; // x=22, y=14
        pixel_data[14][23] = 4'b0000; // x=23, y=14
        pixel_data[14][24] = 4'b0111; // x=24, y=14
        pixel_data[14][25] = 4'b0111; // x=25, y=14
        pixel_data[14][26] = 4'b0111; // x=26, y=14
        pixel_data[14][27] = 4'b0111; // x=27, y=14
        pixel_data[14][28] = 4'b0111; // x=28, y=14
        pixel_data[14][29] = 4'b0111; // x=29, y=14
        pixel_data[14][30] = 4'b0111; // x=30, y=14
        pixel_data[14][31] = 4'b0111; // x=31, y=14
        pixel_data[14][32] = 4'b0111; // x=32, y=14
        pixel_data[14][33] = 4'b0111; // x=33, y=14
        pixel_data[14][34] = 4'b0111; // x=34, y=14
        pixel_data[14][35] = 4'b0111; // x=35, y=14
        pixel_data[14][36] = 4'b0111; // x=36, y=14
        pixel_data[14][37] = 4'b0111; // x=37, y=14
        pixel_data[14][38] = 4'b0111; // x=38, y=14
        pixel_data[14][39] = 4'b0111; // x=39, y=14
        pixel_data[14][40] = 4'b0111; // x=40, y=14
        pixel_data[14][41] = 4'b0111; // x=41, y=14
        pixel_data[14][42] = 4'b0111; // x=42, y=14
        pixel_data[14][43] = 4'b0111; // x=43, y=14
        pixel_data[14][44] = 4'b0111; // x=44, y=14
        pixel_data[14][45] = 4'b0111; // x=45, y=14
        pixel_data[14][46] = 4'b0111; // x=46, y=14
        pixel_data[14][47] = 4'b0111; // x=47, y=14
        pixel_data[14][48] = 4'b0111; // x=48, y=14
        pixel_data[14][49] = 4'b0111; // x=49, y=14
        pixel_data[14][50] = 4'b0111; // x=50, y=14
        pixel_data[14][51] = 4'b0111; // x=51, y=14
        pixel_data[14][52] = 4'b0111; // x=52, y=14
        pixel_data[14][53] = 4'b0111; // x=53, y=14
        pixel_data[14][54] = 4'b0111; // x=54, y=14
        pixel_data[14][55] = 4'b0111; // x=55, y=14
        pixel_data[14][56] = 4'b0111; // x=56, y=14
        pixel_data[14][57] = 4'b0111; // x=57, y=14
        pixel_data[14][58] = 4'b0111; // x=58, y=14
        pixel_data[14][59] = 4'b0111; // x=59, y=14
        pixel_data[14][60] = 4'b0111; // x=60, y=14
        pixel_data[14][61] = 4'b0111; // x=61, y=14
        pixel_data[14][62] = 4'b0111; // x=62, y=14
        pixel_data[14][63] = 4'b0111; // x=63, y=14
        pixel_data[14][64] = 4'b0111; // x=64, y=14
        pixel_data[14][65] = 4'b0111; // x=65, y=14
        pixel_data[14][66] = 4'b0111; // x=66, y=14
        pixel_data[14][67] = 4'b0111; // x=67, y=14
        pixel_data[14][68] = 4'b0111; // x=68, y=14
        pixel_data[14][69] = 4'b0111; // x=69, y=14
        pixel_data[14][70] = 4'b0111; // x=70, y=14
        pixel_data[14][71] = 4'b0111; // x=71, y=14
        pixel_data[14][72] = 4'b0111; // x=72, y=14
        pixel_data[14][73] = 4'b0111; // x=73, y=14
        pixel_data[14][74] = 4'b0111; // x=74, y=14
        pixel_data[14][75] = 4'b0111; // x=75, y=14
        pixel_data[14][76] = 4'b0111; // x=76, y=14
        pixel_data[14][77] = 4'b0111; // x=77, y=14
        pixel_data[14][78] = 4'b0111; // x=78, y=14
        pixel_data[14][79] = 4'b0111; // x=79, y=14
        pixel_data[14][80] = 4'b0111; // x=80, y=14
        pixel_data[14][81] = 4'b0111; // x=81, y=14
        pixel_data[14][82] = 4'b0111; // x=82, y=14
        pixel_data[14][83] = 4'b0111; // x=83, y=14
        pixel_data[14][84] = 4'b0111; // x=84, y=14
        pixel_data[14][85] = 4'b0111; // x=85, y=14
        pixel_data[14][86] = 4'b0111; // x=86, y=14
        pixel_data[14][87] = 4'b0111; // x=87, y=14
        pixel_data[14][88] = 4'b0111; // x=88, y=14
        pixel_data[14][89] = 4'b0111; // x=89, y=14
        pixel_data[14][90] = 4'b0111; // x=90, y=14
        pixel_data[14][91] = 4'b0111; // x=91, y=14
        pixel_data[14][92] = 4'b0111; // x=92, y=14
        pixel_data[14][93] = 4'b0111; // x=93, y=14
        pixel_data[14][94] = 4'b0111; // x=94, y=14
        pixel_data[14][95] = 4'b0111; // x=95, y=14
        pixel_data[14][96] = 4'b0111; // x=96, y=14
        pixel_data[14][97] = 4'b0111; // x=97, y=14
        pixel_data[14][98] = 4'b0111; // x=98, y=14
        pixel_data[14][99] = 4'b0111; // x=99, y=14
        pixel_data[14][100] = 4'b0111; // x=100, y=14
        pixel_data[14][101] = 4'b0111; // x=101, y=14
        pixel_data[14][102] = 4'b0111; // x=102, y=14
        pixel_data[14][103] = 4'b0111; // x=103, y=14
        pixel_data[14][104] = 4'b0111; // x=104, y=14
        pixel_data[14][105] = 4'b0111; // x=105, y=14
        pixel_data[14][106] = 4'b0111; // x=106, y=14
        pixel_data[14][107] = 4'b0111; // x=107, y=14
        pixel_data[14][108] = 4'b0111; // x=108, y=14
        pixel_data[14][109] = 4'b0111; // x=109, y=14
        pixel_data[14][110] = 4'b0111; // x=110, y=14
        pixel_data[14][111] = 4'b0111; // x=111, y=14
        pixel_data[14][112] = 4'b0111; // x=112, y=14
        pixel_data[14][113] = 4'b0111; // x=113, y=14
        pixel_data[14][114] = 4'b0111; // x=114, y=14
        pixel_data[14][115] = 4'b0111; // x=115, y=14
        pixel_data[14][116] = 4'b0111; // x=116, y=14
        pixel_data[14][117] = 4'b0111; // x=117, y=14
        pixel_data[14][118] = 4'b0111; // x=118, y=14
        pixel_data[14][119] = 4'b0111; // x=119, y=14
        pixel_data[14][120] = 4'b0111; // x=120, y=14
        pixel_data[14][121] = 4'b0111; // x=121, y=14
        pixel_data[14][122] = 4'b0111; // x=122, y=14
        pixel_data[14][123] = 4'b0111; // x=123, y=14
        pixel_data[14][124] = 4'b0111; // x=124, y=14
        pixel_data[14][125] = 4'b0111; // x=125, y=14
        pixel_data[14][126] = 4'b0111; // x=126, y=14
        pixel_data[14][127] = 4'b0111; // x=127, y=14
        pixel_data[14][128] = 4'b0111; // x=128, y=14
        pixel_data[14][129] = 4'b0111; // x=129, y=14
        pixel_data[14][130] = 4'b0111; // x=130, y=14
        pixel_data[14][131] = 4'b0111; // x=131, y=14
        pixel_data[14][132] = 4'b0111; // x=132, y=14
        pixel_data[14][133] = 4'b0111; // x=133, y=14
        pixel_data[14][134] = 4'b0111; // x=134, y=14
        pixel_data[14][135] = 4'b0111; // x=135, y=14
        pixel_data[14][136] = 4'b0111; // x=136, y=14
        pixel_data[14][137] = 4'b0111; // x=137, y=14
        pixel_data[14][138] = 4'b0111; // x=138, y=14
        pixel_data[14][139] = 4'b0111; // x=139, y=14
        pixel_data[14][140] = 4'b0111; // x=140, y=14
        pixel_data[14][141] = 4'b0111; // x=141, y=14
        pixel_data[14][142] = 4'b0111; // x=142, y=14
        pixel_data[14][143] = 4'b0111; // x=143, y=14
        pixel_data[14][144] = 4'b0111; // x=144, y=14
        pixel_data[14][145] = 4'b0111; // x=145, y=14
        pixel_data[14][146] = 4'b0111; // x=146, y=14
        pixel_data[14][147] = 4'b0111; // x=147, y=14
        pixel_data[14][148] = 4'b0111; // x=148, y=14
        pixel_data[14][149] = 4'b0111; // x=149, y=14
        pixel_data[14][150] = 4'b0111; // x=150, y=14
        pixel_data[14][151] = 4'b0111; // x=151, y=14
        pixel_data[14][152] = 4'b0111; // x=152, y=14
        pixel_data[14][153] = 4'b0111; // x=153, y=14
        pixel_data[14][154] = 4'b0111; // x=154, y=14
        pixel_data[14][155] = 4'b0111; // x=155, y=14
        pixel_data[14][156] = 4'b0111; // x=156, y=14
        pixel_data[14][157] = 4'b0111; // x=157, y=14
        pixel_data[14][158] = 4'b0111; // x=158, y=14
        pixel_data[14][159] = 4'b0111; // x=159, y=14
        pixel_data[14][160] = 4'b0111; // x=160, y=14
        pixel_data[14][161] = 4'b0111; // x=161, y=14
        pixel_data[14][162] = 4'b0111; // x=162, y=14
        pixel_data[14][163] = 4'b0111; // x=163, y=14
        pixel_data[14][164] = 4'b0111; // x=164, y=14
        pixel_data[14][165] = 4'b0111; // x=165, y=14
        pixel_data[14][166] = 4'b0111; // x=166, y=14
        pixel_data[14][167] = 4'b0111; // x=167, y=14
        pixel_data[14][168] = 4'b0111; // x=168, y=14
        pixel_data[14][169] = 4'b0111; // x=169, y=14
        pixel_data[14][170] = 4'b0111; // x=170, y=14
        pixel_data[14][171] = 4'b0111; // x=171, y=14
        pixel_data[14][172] = 4'b0111; // x=172, y=14
        pixel_data[14][173] = 4'b0111; // x=173, y=14
        pixel_data[14][174] = 4'b0111; // x=174, y=14
        pixel_data[14][175] = 4'b0111; // x=175, y=14
        pixel_data[14][176] = 4'b0111; // x=176, y=14
        pixel_data[14][177] = 4'b0111; // x=177, y=14
        pixel_data[14][178] = 4'b0111; // x=178, y=14
        pixel_data[14][179] = 4'b0111; // x=179, y=14
        pixel_data[15][0] = 4'b0111; // x=0, y=15
        pixel_data[15][1] = 4'b0111; // x=1, y=15
        pixel_data[15][2] = 4'b0111; // x=2, y=15
        pixel_data[15][3] = 4'b0111; // x=3, y=15
        pixel_data[15][4] = 4'b0111; // x=4, y=15
        pixel_data[15][5] = 4'b0111; // x=5, y=15
        pixel_data[15][6] = 4'b0111; // x=6, y=15
        pixel_data[15][7] = 4'b0111; // x=7, y=15
        pixel_data[15][8] = 4'b0111; // x=8, y=15
        pixel_data[15][9] = 4'b0111; // x=9, y=15
        pixel_data[15][10] = 4'b0111; // x=10, y=15
        pixel_data[15][11] = 4'b0111; // x=11, y=15
        pixel_data[15][12] = 4'b0111; // x=12, y=15
        pixel_data[15][13] = 4'b0111; // x=13, y=15
        pixel_data[15][14] = 4'b0111; // x=14, y=15
        pixel_data[15][15] = 4'b0111; // x=15, y=15
        pixel_data[15][16] = 4'b0000; // x=16, y=15
        pixel_data[15][17] = 4'b0000; // x=17, y=15
        pixel_data[15][18] = 4'b0000; // x=18, y=15
        pixel_data[15][19] = 4'b0000; // x=19, y=15
        pixel_data[15][20] = 4'b0111; // x=20, y=15
        pixel_data[15][21] = 4'b0111; // x=21, y=15
        pixel_data[15][22] = 4'b0000; // x=22, y=15
        pixel_data[15][23] = 4'b0000; // x=23, y=15
        pixel_data[15][24] = 4'b0000; // x=24, y=15
        pixel_data[15][25] = 4'b0000; // x=25, y=15
        pixel_data[15][26] = 4'b0000; // x=26, y=15
        pixel_data[15][27] = 4'b0111; // x=27, y=15
        pixel_data[15][28] = 4'b0111; // x=28, y=15
        pixel_data[15][29] = 4'b0111; // x=29, y=15
        pixel_data[15][30] = 4'b0111; // x=30, y=15
        pixel_data[15][31] = 4'b0111; // x=31, y=15
        pixel_data[15][32] = 4'b0111; // x=32, y=15
        pixel_data[15][33] = 4'b0111; // x=33, y=15
        pixel_data[15][34] = 4'b0111; // x=34, y=15
        pixel_data[15][35] = 4'b0111; // x=35, y=15
        pixel_data[15][36] = 4'b0111; // x=36, y=15
        pixel_data[15][37] = 4'b0111; // x=37, y=15
        pixel_data[15][38] = 4'b0111; // x=38, y=15
        pixel_data[15][39] = 4'b0111; // x=39, y=15
        pixel_data[15][40] = 4'b0111; // x=40, y=15
        pixel_data[15][41] = 4'b0111; // x=41, y=15
        pixel_data[15][42] = 4'b0111; // x=42, y=15
        pixel_data[15][43] = 4'b0111; // x=43, y=15
        pixel_data[15][44] = 4'b0111; // x=44, y=15
        pixel_data[15][45] = 4'b0111; // x=45, y=15
        pixel_data[15][46] = 4'b0111; // x=46, y=15
        pixel_data[15][47] = 4'b0111; // x=47, y=15
        pixel_data[15][48] = 4'b0111; // x=48, y=15
        pixel_data[15][49] = 4'b0111; // x=49, y=15
        pixel_data[15][50] = 4'b0111; // x=50, y=15
        pixel_data[15][51] = 4'b0111; // x=51, y=15
        pixel_data[15][52] = 4'b0111; // x=52, y=15
        pixel_data[15][53] = 4'b0111; // x=53, y=15
        pixel_data[15][54] = 4'b0111; // x=54, y=15
        pixel_data[15][55] = 4'b0111; // x=55, y=15
        pixel_data[15][56] = 4'b0111; // x=56, y=15
        pixel_data[15][57] = 4'b0111; // x=57, y=15
        pixel_data[15][58] = 4'b0111; // x=58, y=15
        pixel_data[15][59] = 4'b0111; // x=59, y=15
        pixel_data[15][60] = 4'b0111; // x=60, y=15
        pixel_data[15][61] = 4'b0111; // x=61, y=15
        pixel_data[15][62] = 4'b0111; // x=62, y=15
        pixel_data[15][63] = 4'b0111; // x=63, y=15
        pixel_data[15][64] = 4'b0111; // x=64, y=15
        pixel_data[15][65] = 4'b0111; // x=65, y=15
        pixel_data[15][66] = 4'b0111; // x=66, y=15
        pixel_data[15][67] = 4'b0111; // x=67, y=15
        pixel_data[15][68] = 4'b0111; // x=68, y=15
        pixel_data[15][69] = 4'b0111; // x=69, y=15
        pixel_data[15][70] = 4'b0111; // x=70, y=15
        pixel_data[15][71] = 4'b0111; // x=71, y=15
        pixel_data[15][72] = 4'b0111; // x=72, y=15
        pixel_data[15][73] = 4'b0111; // x=73, y=15
        pixel_data[15][74] = 4'b0111; // x=74, y=15
        pixel_data[15][75] = 4'b0111; // x=75, y=15
        pixel_data[15][76] = 4'b0111; // x=76, y=15
        pixel_data[15][77] = 4'b0111; // x=77, y=15
        pixel_data[15][78] = 4'b0111; // x=78, y=15
        pixel_data[15][79] = 4'b0111; // x=79, y=15
        pixel_data[15][80] = 4'b0111; // x=80, y=15
        pixel_data[15][81] = 4'b0111; // x=81, y=15
        pixel_data[15][82] = 4'b0111; // x=82, y=15
        pixel_data[15][83] = 4'b0111; // x=83, y=15
        pixel_data[15][84] = 4'b0111; // x=84, y=15
        pixel_data[15][85] = 4'b0111; // x=85, y=15
        pixel_data[15][86] = 4'b0111; // x=86, y=15
        pixel_data[15][87] = 4'b0111; // x=87, y=15
        pixel_data[15][88] = 4'b0111; // x=88, y=15
        pixel_data[15][89] = 4'b0111; // x=89, y=15
        pixel_data[15][90] = 4'b0111; // x=90, y=15
        pixel_data[15][91] = 4'b0111; // x=91, y=15
        pixel_data[15][92] = 4'b0111; // x=92, y=15
        pixel_data[15][93] = 4'b0111; // x=93, y=15
        pixel_data[15][94] = 4'b0111; // x=94, y=15
        pixel_data[15][95] = 4'b0111; // x=95, y=15
        pixel_data[15][96] = 4'b0111; // x=96, y=15
        pixel_data[15][97] = 4'b0111; // x=97, y=15
        pixel_data[15][98] = 4'b0111; // x=98, y=15
        pixel_data[15][99] = 4'b0111; // x=99, y=15
        pixel_data[15][100] = 4'b0111; // x=100, y=15
        pixel_data[15][101] = 4'b0111; // x=101, y=15
        pixel_data[15][102] = 4'b0111; // x=102, y=15
        pixel_data[15][103] = 4'b0111; // x=103, y=15
        pixel_data[15][104] = 4'b0111; // x=104, y=15
        pixel_data[15][105] = 4'b0111; // x=105, y=15
        pixel_data[15][106] = 4'b0111; // x=106, y=15
        pixel_data[15][107] = 4'b0111; // x=107, y=15
        pixel_data[15][108] = 4'b0111; // x=108, y=15
        pixel_data[15][109] = 4'b0111; // x=109, y=15
        pixel_data[15][110] = 4'b0111; // x=110, y=15
        pixel_data[15][111] = 4'b0111; // x=111, y=15
        pixel_data[15][112] = 4'b0111; // x=112, y=15
        pixel_data[15][113] = 4'b0111; // x=113, y=15
        pixel_data[15][114] = 4'b0111; // x=114, y=15
        pixel_data[15][115] = 4'b0111; // x=115, y=15
        pixel_data[15][116] = 4'b0111; // x=116, y=15
        pixel_data[15][117] = 4'b0111; // x=117, y=15
        pixel_data[15][118] = 4'b0111; // x=118, y=15
        pixel_data[15][119] = 4'b0111; // x=119, y=15
        pixel_data[15][120] = 4'b0111; // x=120, y=15
        pixel_data[15][121] = 4'b0111; // x=121, y=15
        pixel_data[15][122] = 4'b0111; // x=122, y=15
        pixel_data[15][123] = 4'b0111; // x=123, y=15
        pixel_data[15][124] = 4'b0111; // x=124, y=15
        pixel_data[15][125] = 4'b0111; // x=125, y=15
        pixel_data[15][126] = 4'b0111; // x=126, y=15
        pixel_data[15][127] = 4'b0111; // x=127, y=15
        pixel_data[15][128] = 4'b0111; // x=128, y=15
        pixel_data[15][129] = 4'b0111; // x=129, y=15
        pixel_data[15][130] = 4'b0111; // x=130, y=15
        pixel_data[15][131] = 4'b0111; // x=131, y=15
        pixel_data[15][132] = 4'b0111; // x=132, y=15
        pixel_data[15][133] = 4'b0111; // x=133, y=15
        pixel_data[15][134] = 4'b0111; // x=134, y=15
        pixel_data[15][135] = 4'b0111; // x=135, y=15
        pixel_data[15][136] = 4'b0111; // x=136, y=15
        pixel_data[15][137] = 4'b0111; // x=137, y=15
        pixel_data[15][138] = 4'b0111; // x=138, y=15
        pixel_data[15][139] = 4'b0111; // x=139, y=15
        pixel_data[15][140] = 4'b0111; // x=140, y=15
        pixel_data[15][141] = 4'b0111; // x=141, y=15
        pixel_data[15][142] = 4'b0111; // x=142, y=15
        pixel_data[15][143] = 4'b0111; // x=143, y=15
        pixel_data[15][144] = 4'b0111; // x=144, y=15
        pixel_data[15][145] = 4'b0111; // x=145, y=15
        pixel_data[15][146] = 4'b0111; // x=146, y=15
        pixel_data[15][147] = 4'b0111; // x=147, y=15
        pixel_data[15][148] = 4'b0111; // x=148, y=15
        pixel_data[15][149] = 4'b0111; // x=149, y=15
        pixel_data[15][150] = 4'b0111; // x=150, y=15
        pixel_data[15][151] = 4'b0111; // x=151, y=15
        pixel_data[15][152] = 4'b0111; // x=152, y=15
        pixel_data[15][153] = 4'b0111; // x=153, y=15
        pixel_data[15][154] = 4'b0111; // x=154, y=15
        pixel_data[15][155] = 4'b0111; // x=155, y=15
        pixel_data[15][156] = 4'b0111; // x=156, y=15
        pixel_data[15][157] = 4'b0111; // x=157, y=15
        pixel_data[15][158] = 4'b0111; // x=158, y=15
        pixel_data[15][159] = 4'b0111; // x=159, y=15
        pixel_data[15][160] = 4'b0111; // x=160, y=15
        pixel_data[15][161] = 4'b0111; // x=161, y=15
        pixel_data[15][162] = 4'b0111; // x=162, y=15
        pixel_data[15][163] = 4'b0111; // x=163, y=15
        pixel_data[15][164] = 4'b0111; // x=164, y=15
        pixel_data[15][165] = 4'b0111; // x=165, y=15
        pixel_data[15][166] = 4'b0111; // x=166, y=15
        pixel_data[15][167] = 4'b0111; // x=167, y=15
        pixel_data[15][168] = 4'b0111; // x=168, y=15
        pixel_data[15][169] = 4'b0111; // x=169, y=15
        pixel_data[15][170] = 4'b0111; // x=170, y=15
        pixel_data[15][171] = 4'b0111; // x=171, y=15
        pixel_data[15][172] = 4'b0111; // x=172, y=15
        pixel_data[15][173] = 4'b0111; // x=173, y=15
        pixel_data[15][174] = 4'b0111; // x=174, y=15
        pixel_data[15][175] = 4'b0111; // x=175, y=15
        pixel_data[15][176] = 4'b0111; // x=176, y=15
        pixel_data[15][177] = 4'b0111; // x=177, y=15
        pixel_data[15][178] = 4'b0111; // x=178, y=15
        pixel_data[15][179] = 4'b0111; // x=179, y=15
        pixel_data[16][0] = 4'b0111; // x=0, y=16
        pixel_data[16][1] = 4'b0111; // x=1, y=16
        pixel_data[16][2] = 4'b0111; // x=2, y=16
        pixel_data[16][3] = 4'b0111; // x=3, y=16
        pixel_data[16][4] = 4'b0111; // x=4, y=16
        pixel_data[16][5] = 4'b0111; // x=5, y=16
        pixel_data[16][6] = 4'b0111; // x=6, y=16
        pixel_data[16][7] = 4'b0111; // x=7, y=16
        pixel_data[16][8] = 4'b0111; // x=8, y=16
        pixel_data[16][9] = 4'b0111; // x=9, y=16
        pixel_data[16][10] = 4'b0111; // x=10, y=16
        pixel_data[16][11] = 4'b0111; // x=11, y=16
        pixel_data[16][12] = 4'b0111; // x=12, y=16
        pixel_data[16][13] = 4'b0111; // x=13, y=16
        pixel_data[16][14] = 4'b0000; // x=14, y=16
        pixel_data[16][15] = 4'b0111; // x=15, y=16
        pixel_data[16][16] = 4'b0111; // x=16, y=16
        pixel_data[16][17] = 4'b0111; // x=17, y=16
        pixel_data[16][18] = 4'b0111; // x=18, y=16
        pixel_data[16][19] = 4'b0111; // x=19, y=16
        pixel_data[16][20] = 4'b0111; // x=20, y=16
        pixel_data[16][21] = 4'b0111; // x=21, y=16
        pixel_data[16][22] = 4'b0111; // x=22, y=16
        pixel_data[16][23] = 4'b0111; // x=23, y=16
        pixel_data[16][24] = 4'b0111; // x=24, y=16
        pixel_data[16][25] = 4'b0111; // x=25, y=16
        pixel_data[16][26] = 4'b0111; // x=26, y=16
        pixel_data[16][27] = 4'b0111; // x=27, y=16
        pixel_data[16][28] = 4'b0111; // x=28, y=16
        pixel_data[16][29] = 4'b0111; // x=29, y=16
        pixel_data[16][30] = 4'b0111; // x=30, y=16
        pixel_data[16][31] = 4'b0111; // x=31, y=16
        pixel_data[16][32] = 4'b0111; // x=32, y=16
        pixel_data[16][33] = 4'b0111; // x=33, y=16
        pixel_data[16][34] = 4'b0111; // x=34, y=16
        pixel_data[16][35] = 4'b0111; // x=35, y=16
        pixel_data[16][36] = 4'b0111; // x=36, y=16
        pixel_data[16][37] = 4'b0111; // x=37, y=16
        pixel_data[16][38] = 4'b0111; // x=38, y=16
        pixel_data[16][39] = 4'b0111; // x=39, y=16
        pixel_data[16][40] = 4'b0111; // x=40, y=16
        pixel_data[16][41] = 4'b0111; // x=41, y=16
        pixel_data[16][42] = 4'b0111; // x=42, y=16
        pixel_data[16][43] = 4'b0111; // x=43, y=16
        pixel_data[16][44] = 4'b0111; // x=44, y=16
        pixel_data[16][45] = 4'b0111; // x=45, y=16
        pixel_data[16][46] = 4'b0111; // x=46, y=16
        pixel_data[16][47] = 4'b0111; // x=47, y=16
        pixel_data[16][48] = 4'b0111; // x=48, y=16
        pixel_data[16][49] = 4'b0111; // x=49, y=16
        pixel_data[16][50] = 4'b0111; // x=50, y=16
        pixel_data[16][51] = 4'b0111; // x=51, y=16
        pixel_data[16][52] = 4'b0111; // x=52, y=16
        pixel_data[16][53] = 4'b0111; // x=53, y=16
        pixel_data[16][54] = 4'b0111; // x=54, y=16
        pixel_data[16][55] = 4'b0111; // x=55, y=16
        pixel_data[16][56] = 4'b0111; // x=56, y=16
        pixel_data[16][57] = 4'b0111; // x=57, y=16
        pixel_data[16][58] = 4'b0111; // x=58, y=16
        pixel_data[16][59] = 4'b0111; // x=59, y=16
        pixel_data[16][60] = 4'b0111; // x=60, y=16
        pixel_data[16][61] = 4'b0111; // x=61, y=16
        pixel_data[16][62] = 4'b0111; // x=62, y=16
        pixel_data[16][63] = 4'b0111; // x=63, y=16
        pixel_data[16][64] = 4'b0111; // x=64, y=16
        pixel_data[16][65] = 4'b0111; // x=65, y=16
        pixel_data[16][66] = 4'b0111; // x=66, y=16
        pixel_data[16][67] = 4'b0111; // x=67, y=16
        pixel_data[16][68] = 4'b0111; // x=68, y=16
        pixel_data[16][69] = 4'b0111; // x=69, y=16
        pixel_data[16][70] = 4'b0111; // x=70, y=16
        pixel_data[16][71] = 4'b0111; // x=71, y=16
        pixel_data[16][72] = 4'b0111; // x=72, y=16
        pixel_data[16][73] = 4'b0111; // x=73, y=16
        pixel_data[16][74] = 4'b0111; // x=74, y=16
        pixel_data[16][75] = 4'b0111; // x=75, y=16
        pixel_data[16][76] = 4'b0111; // x=76, y=16
        pixel_data[16][77] = 4'b0111; // x=77, y=16
        pixel_data[16][78] = 4'b0111; // x=78, y=16
        pixel_data[16][79] = 4'b0111; // x=79, y=16
        pixel_data[16][80] = 4'b0111; // x=80, y=16
        pixel_data[16][81] = 4'b0111; // x=81, y=16
        pixel_data[16][82] = 4'b0111; // x=82, y=16
        pixel_data[16][83] = 4'b0111; // x=83, y=16
        pixel_data[16][84] = 4'b0111; // x=84, y=16
        pixel_data[16][85] = 4'b0111; // x=85, y=16
        pixel_data[16][86] = 4'b0111; // x=86, y=16
        pixel_data[16][87] = 4'b0111; // x=87, y=16
        pixel_data[16][88] = 4'b0111; // x=88, y=16
        pixel_data[16][89] = 4'b0111; // x=89, y=16
        pixel_data[16][90] = 4'b0111; // x=90, y=16
        pixel_data[16][91] = 4'b0111; // x=91, y=16
        pixel_data[16][92] = 4'b0111; // x=92, y=16
        pixel_data[16][93] = 4'b0111; // x=93, y=16
        pixel_data[16][94] = 4'b0111; // x=94, y=16
        pixel_data[16][95] = 4'b0111; // x=95, y=16
        pixel_data[16][96] = 4'b0111; // x=96, y=16
        pixel_data[16][97] = 4'b0111; // x=97, y=16
        pixel_data[16][98] = 4'b0111; // x=98, y=16
        pixel_data[16][99] = 4'b0111; // x=99, y=16
        pixel_data[16][100] = 4'b0111; // x=100, y=16
        pixel_data[16][101] = 4'b0111; // x=101, y=16
        pixel_data[16][102] = 4'b0111; // x=102, y=16
        pixel_data[16][103] = 4'b0111; // x=103, y=16
        pixel_data[16][104] = 4'b0111; // x=104, y=16
        pixel_data[16][105] = 4'b0111; // x=105, y=16
        pixel_data[16][106] = 4'b0111; // x=106, y=16
        pixel_data[16][107] = 4'b0111; // x=107, y=16
        pixel_data[16][108] = 4'b0111; // x=108, y=16
        pixel_data[16][109] = 4'b0111; // x=109, y=16
        pixel_data[16][110] = 4'b0111; // x=110, y=16
        pixel_data[16][111] = 4'b0111; // x=111, y=16
        pixel_data[16][112] = 4'b0111; // x=112, y=16
        pixel_data[16][113] = 4'b0111; // x=113, y=16
        pixel_data[16][114] = 4'b0111; // x=114, y=16
        pixel_data[16][115] = 4'b0111; // x=115, y=16
        pixel_data[16][116] = 4'b0111; // x=116, y=16
        pixel_data[16][117] = 4'b0111; // x=117, y=16
        pixel_data[16][118] = 4'b0111; // x=118, y=16
        pixel_data[16][119] = 4'b0111; // x=119, y=16
        pixel_data[16][120] = 4'b0111; // x=120, y=16
        pixel_data[16][121] = 4'b0111; // x=121, y=16
        pixel_data[16][122] = 4'b0111; // x=122, y=16
        pixel_data[16][123] = 4'b0111; // x=123, y=16
        pixel_data[16][124] = 4'b0111; // x=124, y=16
        pixel_data[16][125] = 4'b0111; // x=125, y=16
        pixel_data[16][126] = 4'b0111; // x=126, y=16
        pixel_data[16][127] = 4'b0111; // x=127, y=16
        pixel_data[16][128] = 4'b0111; // x=128, y=16
        pixel_data[16][129] = 4'b0111; // x=129, y=16
        pixel_data[16][130] = 4'b0111; // x=130, y=16
        pixel_data[16][131] = 4'b0111; // x=131, y=16
        pixel_data[16][132] = 4'b0111; // x=132, y=16
        pixel_data[16][133] = 4'b0111; // x=133, y=16
        pixel_data[16][134] = 4'b0111; // x=134, y=16
        pixel_data[16][135] = 4'b0111; // x=135, y=16
        pixel_data[16][136] = 4'b0111; // x=136, y=16
        pixel_data[16][137] = 4'b0111; // x=137, y=16
        pixel_data[16][138] = 4'b0111; // x=138, y=16
        pixel_data[16][139] = 4'b0111; // x=139, y=16
        pixel_data[16][140] = 4'b0111; // x=140, y=16
        pixel_data[16][141] = 4'b0111; // x=141, y=16
        pixel_data[16][142] = 4'b0111; // x=142, y=16
        pixel_data[16][143] = 4'b0111; // x=143, y=16
        pixel_data[16][144] = 4'b0111; // x=144, y=16
        pixel_data[16][145] = 4'b0111; // x=145, y=16
        pixel_data[16][146] = 4'b0111; // x=146, y=16
        pixel_data[16][147] = 4'b0111; // x=147, y=16
        pixel_data[16][148] = 4'b0111; // x=148, y=16
        pixel_data[16][149] = 4'b0111; // x=149, y=16
        pixel_data[16][150] = 4'b0111; // x=150, y=16
        pixel_data[16][151] = 4'b0111; // x=151, y=16
        pixel_data[16][152] = 4'b0111; // x=152, y=16
        pixel_data[16][153] = 4'b0111; // x=153, y=16
        pixel_data[16][154] = 4'b0111; // x=154, y=16
        pixel_data[16][155] = 4'b0111; // x=155, y=16
        pixel_data[16][156] = 4'b0111; // x=156, y=16
        pixel_data[16][157] = 4'b0111; // x=157, y=16
        pixel_data[16][158] = 4'b0111; // x=158, y=16
        pixel_data[16][159] = 4'b0111; // x=159, y=16
        pixel_data[16][160] = 4'b0111; // x=160, y=16
        pixel_data[16][161] = 4'b0111; // x=161, y=16
        pixel_data[16][162] = 4'b0111; // x=162, y=16
        pixel_data[16][163] = 4'b0111; // x=163, y=16
        pixel_data[16][164] = 4'b0111; // x=164, y=16
        pixel_data[16][165] = 4'b0111; // x=165, y=16
        pixel_data[16][166] = 4'b0111; // x=166, y=16
        pixel_data[16][167] = 4'b0111; // x=167, y=16
        pixel_data[16][168] = 4'b0111; // x=168, y=16
        pixel_data[16][169] = 4'b0111; // x=169, y=16
        pixel_data[16][170] = 4'b0111; // x=170, y=16
        pixel_data[16][171] = 4'b0111; // x=171, y=16
        pixel_data[16][172] = 4'b0111; // x=172, y=16
        pixel_data[16][173] = 4'b0111; // x=173, y=16
        pixel_data[16][174] = 4'b0111; // x=174, y=16
        pixel_data[16][175] = 4'b0111; // x=175, y=16
        pixel_data[16][176] = 4'b0111; // x=176, y=16
        pixel_data[16][177] = 4'b0111; // x=177, y=16
        pixel_data[16][178] = 4'b0111; // x=178, y=16
        pixel_data[16][179] = 4'b0111; // x=179, y=16
        pixel_data[17][0] = 4'b0111; // x=0, y=17
        pixel_data[17][1] = 4'b0111; // x=1, y=17
        pixel_data[17][2] = 4'b0111; // x=2, y=17
        pixel_data[17][3] = 4'b0111; // x=3, y=17
        pixel_data[17][4] = 4'b0111; // x=4, y=17
        pixel_data[17][5] = 4'b0111; // x=5, y=17
        pixel_data[17][6] = 4'b0111; // x=6, y=17
        pixel_data[17][7] = 4'b0111; // x=7, y=17
        pixel_data[17][8] = 4'b0111; // x=8, y=17
        pixel_data[17][9] = 4'b0111; // x=9, y=17
        pixel_data[17][10] = 4'b0111; // x=10, y=17
        pixel_data[17][11] = 4'b0111; // x=11, y=17
        pixel_data[17][12] = 4'b0000; // x=12, y=17
        pixel_data[17][13] = 4'b0111; // x=13, y=17
        pixel_data[17][14] = 4'b0111; // x=14, y=17
        pixel_data[17][15] = 4'b1110; // x=15, y=17
        pixel_data[17][16] = 4'b1001; // x=16, y=17
        pixel_data[17][17] = 4'b0010; // x=17, y=17
        pixel_data[17][18] = 4'b1000; // x=18, y=17
        pixel_data[17][19] = 4'b1100; // x=19, y=17
        pixel_data[17][20] = 4'b0011; // x=20, y=17
        pixel_data[17][21] = 4'b0011; // x=21, y=17
        pixel_data[17][22] = 4'b1100; // x=22, y=17
        pixel_data[17][23] = 4'b1000; // x=23, y=17
        pixel_data[17][24] = 4'b0101; // x=24, y=17
        pixel_data[17][25] = 4'b1001; // x=25, y=17
        pixel_data[17][26] = 4'b1110; // x=26, y=17
        pixel_data[17][27] = 4'b0111; // x=27, y=17
        pixel_data[17][28] = 4'b0111; // x=28, y=17
        pixel_data[17][29] = 4'b0000; // x=29, y=17
        pixel_data[17][30] = 4'b0111; // x=30, y=17
        pixel_data[17][31] = 4'b0111; // x=31, y=17
        pixel_data[17][32] = 4'b0111; // x=32, y=17
        pixel_data[17][33] = 4'b0111; // x=33, y=17
        pixel_data[17][34] = 4'b0111; // x=34, y=17
        pixel_data[17][35] = 4'b0111; // x=35, y=17
        pixel_data[17][36] = 4'b0111; // x=36, y=17
        pixel_data[17][37] = 4'b0111; // x=37, y=17
        pixel_data[17][38] = 4'b0111; // x=38, y=17
        pixel_data[17][39] = 4'b0111; // x=39, y=17
        pixel_data[17][40] = 4'b0111; // x=40, y=17
        pixel_data[17][41] = 4'b0111; // x=41, y=17
        pixel_data[17][42] = 4'b0111; // x=42, y=17
        pixel_data[17][43] = 4'b0111; // x=43, y=17
        pixel_data[17][44] = 4'b0111; // x=44, y=17
        pixel_data[17][45] = 4'b0111; // x=45, y=17
        pixel_data[17][46] = 4'b0111; // x=46, y=17
        pixel_data[17][47] = 4'b0111; // x=47, y=17
        pixel_data[17][48] = 4'b0111; // x=48, y=17
        pixel_data[17][49] = 4'b0111; // x=49, y=17
        pixel_data[17][50] = 4'b0111; // x=50, y=17
        pixel_data[17][51] = 4'b0111; // x=51, y=17
        pixel_data[17][52] = 4'b0111; // x=52, y=17
        pixel_data[17][53] = 4'b0111; // x=53, y=17
        pixel_data[17][54] = 4'b0111; // x=54, y=17
        pixel_data[17][55] = 4'b0111; // x=55, y=17
        pixel_data[17][56] = 4'b0111; // x=56, y=17
        pixel_data[17][57] = 4'b0111; // x=57, y=17
        pixel_data[17][58] = 4'b0111; // x=58, y=17
        pixel_data[17][59] = 4'b0111; // x=59, y=17
        pixel_data[17][60] = 4'b0111; // x=60, y=17
        pixel_data[17][61] = 4'b0111; // x=61, y=17
        pixel_data[17][62] = 4'b0111; // x=62, y=17
        pixel_data[17][63] = 4'b0111; // x=63, y=17
        pixel_data[17][64] = 4'b0111; // x=64, y=17
        pixel_data[17][65] = 4'b0111; // x=65, y=17
        pixel_data[17][66] = 4'b0111; // x=66, y=17
        pixel_data[17][67] = 4'b0111; // x=67, y=17
        pixel_data[17][68] = 4'b0111; // x=68, y=17
        pixel_data[17][69] = 4'b0111; // x=69, y=17
        pixel_data[17][70] = 4'b0111; // x=70, y=17
        pixel_data[17][71] = 4'b0111; // x=71, y=17
        pixel_data[17][72] = 4'b0111; // x=72, y=17
        pixel_data[17][73] = 4'b0111; // x=73, y=17
        pixel_data[17][74] = 4'b0111; // x=74, y=17
        pixel_data[17][75] = 4'b0111; // x=75, y=17
        pixel_data[17][76] = 4'b0111; // x=76, y=17
        pixel_data[17][77] = 4'b0111; // x=77, y=17
        pixel_data[17][78] = 4'b0111; // x=78, y=17
        pixel_data[17][79] = 4'b0111; // x=79, y=17
        pixel_data[17][80] = 4'b0111; // x=80, y=17
        pixel_data[17][81] = 4'b0111; // x=81, y=17
        pixel_data[17][82] = 4'b0111; // x=82, y=17
        pixel_data[17][83] = 4'b0111; // x=83, y=17
        pixel_data[17][84] = 4'b0111; // x=84, y=17
        pixel_data[17][85] = 4'b0111; // x=85, y=17
        pixel_data[17][86] = 4'b0111; // x=86, y=17
        pixel_data[17][87] = 4'b0111; // x=87, y=17
        pixel_data[17][88] = 4'b0111; // x=88, y=17
        pixel_data[17][89] = 4'b0111; // x=89, y=17
        pixel_data[17][90] = 4'b0111; // x=90, y=17
        pixel_data[17][91] = 4'b0111; // x=91, y=17
        pixel_data[17][92] = 4'b0111; // x=92, y=17
        pixel_data[17][93] = 4'b0111; // x=93, y=17
        pixel_data[17][94] = 4'b0111; // x=94, y=17
        pixel_data[17][95] = 4'b0111; // x=95, y=17
        pixel_data[17][96] = 4'b0111; // x=96, y=17
        pixel_data[17][97] = 4'b0111; // x=97, y=17
        pixel_data[17][98] = 4'b0111; // x=98, y=17
        pixel_data[17][99] = 4'b0111; // x=99, y=17
        pixel_data[17][100] = 4'b0111; // x=100, y=17
        pixel_data[17][101] = 4'b0111; // x=101, y=17
        pixel_data[17][102] = 4'b0111; // x=102, y=17
        pixel_data[17][103] = 4'b0111; // x=103, y=17
        pixel_data[17][104] = 4'b0111; // x=104, y=17
        pixel_data[17][105] = 4'b0111; // x=105, y=17
        pixel_data[17][106] = 4'b0111; // x=106, y=17
        pixel_data[17][107] = 4'b0111; // x=107, y=17
        pixel_data[17][108] = 4'b0111; // x=108, y=17
        pixel_data[17][109] = 4'b0111; // x=109, y=17
        pixel_data[17][110] = 4'b0111; // x=110, y=17
        pixel_data[17][111] = 4'b0111; // x=111, y=17
        pixel_data[17][112] = 4'b0111; // x=112, y=17
        pixel_data[17][113] = 4'b0111; // x=113, y=17
        pixel_data[17][114] = 4'b0111; // x=114, y=17
        pixel_data[17][115] = 4'b0111; // x=115, y=17
        pixel_data[17][116] = 4'b0111; // x=116, y=17
        pixel_data[17][117] = 4'b0111; // x=117, y=17
        pixel_data[17][118] = 4'b0111; // x=118, y=17
        pixel_data[17][119] = 4'b0111; // x=119, y=17
        pixel_data[17][120] = 4'b0111; // x=120, y=17
        pixel_data[17][121] = 4'b0111; // x=121, y=17
        pixel_data[17][122] = 4'b0111; // x=122, y=17
        pixel_data[17][123] = 4'b0111; // x=123, y=17
        pixel_data[17][124] = 4'b0111; // x=124, y=17
        pixel_data[17][125] = 4'b0111; // x=125, y=17
        pixel_data[17][126] = 4'b0111; // x=126, y=17
        pixel_data[17][127] = 4'b0111; // x=127, y=17
        pixel_data[17][128] = 4'b0111; // x=128, y=17
        pixel_data[17][129] = 4'b0111; // x=129, y=17
        pixel_data[17][130] = 4'b0111; // x=130, y=17
        pixel_data[17][131] = 4'b0111; // x=131, y=17
        pixel_data[17][132] = 4'b0111; // x=132, y=17
        pixel_data[17][133] = 4'b0111; // x=133, y=17
        pixel_data[17][134] = 4'b0111; // x=134, y=17
        pixel_data[17][135] = 4'b0111; // x=135, y=17
        pixel_data[17][136] = 4'b0111; // x=136, y=17
        pixel_data[17][137] = 4'b0111; // x=137, y=17
        pixel_data[17][138] = 4'b0111; // x=138, y=17
        pixel_data[17][139] = 4'b0111; // x=139, y=17
        pixel_data[17][140] = 4'b0111; // x=140, y=17
        pixel_data[17][141] = 4'b0111; // x=141, y=17
        pixel_data[17][142] = 4'b0111; // x=142, y=17
        pixel_data[17][143] = 4'b0111; // x=143, y=17
        pixel_data[17][144] = 4'b0111; // x=144, y=17
        pixel_data[17][145] = 4'b0111; // x=145, y=17
        pixel_data[17][146] = 4'b0111; // x=146, y=17
        pixel_data[17][147] = 4'b0111; // x=147, y=17
        pixel_data[17][148] = 4'b0111; // x=148, y=17
        pixel_data[17][149] = 4'b0111; // x=149, y=17
        pixel_data[17][150] = 4'b0111; // x=150, y=17
        pixel_data[17][151] = 4'b0111; // x=151, y=17
        pixel_data[17][152] = 4'b0111; // x=152, y=17
        pixel_data[17][153] = 4'b0111; // x=153, y=17
        pixel_data[17][154] = 4'b0111; // x=154, y=17
        pixel_data[17][155] = 4'b0111; // x=155, y=17
        pixel_data[17][156] = 4'b0111; // x=156, y=17
        pixel_data[17][157] = 4'b0111; // x=157, y=17
        pixel_data[17][158] = 4'b0111; // x=158, y=17
        pixel_data[17][159] = 4'b0111; // x=159, y=17
        pixel_data[17][160] = 4'b0111; // x=160, y=17
        pixel_data[17][161] = 4'b0111; // x=161, y=17
        pixel_data[17][162] = 4'b0111; // x=162, y=17
        pixel_data[17][163] = 4'b0111; // x=163, y=17
        pixel_data[17][164] = 4'b0111; // x=164, y=17
        pixel_data[17][165] = 4'b0111; // x=165, y=17
        pixel_data[17][166] = 4'b0111; // x=166, y=17
        pixel_data[17][167] = 4'b0111; // x=167, y=17
        pixel_data[17][168] = 4'b0111; // x=168, y=17
        pixel_data[17][169] = 4'b0111; // x=169, y=17
        pixel_data[17][170] = 4'b0111; // x=170, y=17
        pixel_data[17][171] = 4'b0111; // x=171, y=17
        pixel_data[17][172] = 4'b0111; // x=172, y=17
        pixel_data[17][173] = 4'b0111; // x=173, y=17
        pixel_data[17][174] = 4'b0111; // x=174, y=17
        pixel_data[17][175] = 4'b0111; // x=175, y=17
        pixel_data[17][176] = 4'b0111; // x=176, y=17
        pixel_data[17][177] = 4'b0111; // x=177, y=17
        pixel_data[17][178] = 4'b0111; // x=178, y=17
        pixel_data[17][179] = 4'b0111; // x=179, y=17
        pixel_data[18][0] = 4'b0111; // x=0, y=18
        pixel_data[18][1] = 4'b0111; // x=1, y=18
        pixel_data[18][2] = 4'b0111; // x=2, y=18
        pixel_data[18][3] = 4'b0111; // x=3, y=18
        pixel_data[18][4] = 4'b0111; // x=4, y=18
        pixel_data[18][5] = 4'b0111; // x=5, y=18
        pixel_data[18][6] = 4'b0111; // x=6, y=18
        pixel_data[18][7] = 4'b0111; // x=7, y=18
        pixel_data[18][8] = 4'b0111; // x=8, y=18
        pixel_data[18][9] = 4'b0111; // x=9, y=18
        pixel_data[18][10] = 4'b0000; // x=10, y=18
        pixel_data[18][11] = 4'b0000; // x=11, y=18
        pixel_data[18][12] = 4'b0111; // x=12, y=18
        pixel_data[18][13] = 4'b0110; // x=13, y=18
        pixel_data[18][14] = 4'b0101; // x=14, y=18
        pixel_data[18][15] = 4'b1011; // x=15, y=18
        pixel_data[18][16] = 4'b1101; // x=16, y=18
        pixel_data[18][17] = 4'b1101; // x=17, y=18
        pixel_data[18][18] = 4'b1101; // x=18, y=18
        pixel_data[18][19] = 4'b1101; // x=19, y=18
        pixel_data[18][20] = 4'b1101; // x=20, y=18
        pixel_data[18][21] = 4'b1101; // x=21, y=18
        pixel_data[18][22] = 4'b1101; // x=22, y=18
        pixel_data[18][23] = 4'b1101; // x=23, y=18
        pixel_data[18][24] = 4'b1101; // x=24, y=18
        pixel_data[18][25] = 4'b1101; // x=25, y=18
        pixel_data[18][26] = 4'b1011; // x=26, y=18
        pixel_data[18][27] = 4'b1000; // x=27, y=18
        pixel_data[18][28] = 4'b0100; // x=28, y=18
        pixel_data[18][29] = 4'b0111; // x=29, y=18
        pixel_data[18][30] = 4'b0000; // x=30, y=18
        pixel_data[18][31] = 4'b0000; // x=31, y=18
        pixel_data[18][32] = 4'b0111; // x=32, y=18
        pixel_data[18][33] = 4'b0111; // x=33, y=18
        pixel_data[18][34] = 4'b0111; // x=34, y=18
        pixel_data[18][35] = 4'b0111; // x=35, y=18
        pixel_data[18][36] = 4'b0111; // x=36, y=18
        pixel_data[18][37] = 4'b0111; // x=37, y=18
        pixel_data[18][38] = 4'b0111; // x=38, y=18
        pixel_data[18][39] = 4'b0111; // x=39, y=18
        pixel_data[18][40] = 4'b0111; // x=40, y=18
        pixel_data[18][41] = 4'b0111; // x=41, y=18
        pixel_data[18][42] = 4'b0111; // x=42, y=18
        pixel_data[18][43] = 4'b0111; // x=43, y=18
        pixel_data[18][44] = 4'b0111; // x=44, y=18
        pixel_data[18][45] = 4'b0111; // x=45, y=18
        pixel_data[18][46] = 4'b0111; // x=46, y=18
        pixel_data[18][47] = 4'b0111; // x=47, y=18
        pixel_data[18][48] = 4'b0111; // x=48, y=18
        pixel_data[18][49] = 4'b0111; // x=49, y=18
        pixel_data[18][50] = 4'b0111; // x=50, y=18
        pixel_data[18][51] = 4'b0111; // x=51, y=18
        pixel_data[18][52] = 4'b0111; // x=52, y=18
        pixel_data[18][53] = 4'b0111; // x=53, y=18
        pixel_data[18][54] = 4'b0111; // x=54, y=18
        pixel_data[18][55] = 4'b0111; // x=55, y=18
        pixel_data[18][56] = 4'b0111; // x=56, y=18
        pixel_data[18][57] = 4'b0111; // x=57, y=18
        pixel_data[18][58] = 4'b0111; // x=58, y=18
        pixel_data[18][59] = 4'b0111; // x=59, y=18
        pixel_data[18][60] = 4'b0111; // x=60, y=18
        pixel_data[18][61] = 4'b0111; // x=61, y=18
        pixel_data[18][62] = 4'b0111; // x=62, y=18
        pixel_data[18][63] = 4'b0111; // x=63, y=18
        pixel_data[18][64] = 4'b0111; // x=64, y=18
        pixel_data[18][65] = 4'b0111; // x=65, y=18
        pixel_data[18][66] = 4'b0111; // x=66, y=18
        pixel_data[18][67] = 4'b0111; // x=67, y=18
        pixel_data[18][68] = 4'b0111; // x=68, y=18
        pixel_data[18][69] = 4'b0111; // x=69, y=18
        pixel_data[18][70] = 4'b0111; // x=70, y=18
        pixel_data[18][71] = 4'b0111; // x=71, y=18
        pixel_data[18][72] = 4'b0111; // x=72, y=18
        pixel_data[18][73] = 4'b0111; // x=73, y=18
        pixel_data[18][74] = 4'b0111; // x=74, y=18
        pixel_data[18][75] = 4'b0111; // x=75, y=18
        pixel_data[18][76] = 4'b0111; // x=76, y=18
        pixel_data[18][77] = 4'b0111; // x=77, y=18
        pixel_data[18][78] = 4'b0111; // x=78, y=18
        pixel_data[18][79] = 4'b0111; // x=79, y=18
        pixel_data[18][80] = 4'b0111; // x=80, y=18
        pixel_data[18][81] = 4'b0111; // x=81, y=18
        pixel_data[18][82] = 4'b0111; // x=82, y=18
        pixel_data[18][83] = 4'b0111; // x=83, y=18
        pixel_data[18][84] = 4'b0111; // x=84, y=18
        pixel_data[18][85] = 4'b0111; // x=85, y=18
        pixel_data[18][86] = 4'b0111; // x=86, y=18
        pixel_data[18][87] = 4'b0111; // x=87, y=18
        pixel_data[18][88] = 4'b0111; // x=88, y=18
        pixel_data[18][89] = 4'b0111; // x=89, y=18
        pixel_data[18][90] = 4'b0111; // x=90, y=18
        pixel_data[18][91] = 4'b0111; // x=91, y=18
        pixel_data[18][92] = 4'b0111; // x=92, y=18
        pixel_data[18][93] = 4'b0111; // x=93, y=18
        pixel_data[18][94] = 4'b0111; // x=94, y=18
        pixel_data[18][95] = 4'b0111; // x=95, y=18
        pixel_data[18][96] = 4'b0111; // x=96, y=18
        pixel_data[18][97] = 4'b0111; // x=97, y=18
        pixel_data[18][98] = 4'b0111; // x=98, y=18
        pixel_data[18][99] = 4'b0111; // x=99, y=18
        pixel_data[18][100] = 4'b0111; // x=100, y=18
        pixel_data[18][101] = 4'b0111; // x=101, y=18
        pixel_data[18][102] = 4'b0111; // x=102, y=18
        pixel_data[18][103] = 4'b0111; // x=103, y=18
        pixel_data[18][104] = 4'b0111; // x=104, y=18
        pixel_data[18][105] = 4'b0111; // x=105, y=18
        pixel_data[18][106] = 4'b0111; // x=106, y=18
        pixel_data[18][107] = 4'b0111; // x=107, y=18
        pixel_data[18][108] = 4'b0111; // x=108, y=18
        pixel_data[18][109] = 4'b0111; // x=109, y=18
        pixel_data[18][110] = 4'b0111; // x=110, y=18
        pixel_data[18][111] = 4'b0111; // x=111, y=18
        pixel_data[18][112] = 4'b0111; // x=112, y=18
        pixel_data[18][113] = 4'b0111; // x=113, y=18
        pixel_data[18][114] = 4'b0111; // x=114, y=18
        pixel_data[18][115] = 4'b0111; // x=115, y=18
        pixel_data[18][116] = 4'b0111; // x=116, y=18
        pixel_data[18][117] = 4'b0111; // x=117, y=18
        pixel_data[18][118] = 4'b0111; // x=118, y=18
        pixel_data[18][119] = 4'b0111; // x=119, y=18
        pixel_data[18][120] = 4'b0111; // x=120, y=18
        pixel_data[18][121] = 4'b0111; // x=121, y=18
        pixel_data[18][122] = 4'b0111; // x=122, y=18
        pixel_data[18][123] = 4'b0111; // x=123, y=18
        pixel_data[18][124] = 4'b0111; // x=124, y=18
        pixel_data[18][125] = 4'b0111; // x=125, y=18
        pixel_data[18][126] = 4'b0111; // x=126, y=18
        pixel_data[18][127] = 4'b0111; // x=127, y=18
        pixel_data[18][128] = 4'b0111; // x=128, y=18
        pixel_data[18][129] = 4'b0111; // x=129, y=18
        pixel_data[18][130] = 4'b0111; // x=130, y=18
        pixel_data[18][131] = 4'b0111; // x=131, y=18
        pixel_data[18][132] = 4'b0111; // x=132, y=18
        pixel_data[18][133] = 4'b0111; // x=133, y=18
        pixel_data[18][134] = 4'b0111; // x=134, y=18
        pixel_data[18][135] = 4'b0111; // x=135, y=18
        pixel_data[18][136] = 4'b0111; // x=136, y=18
        pixel_data[18][137] = 4'b0111; // x=137, y=18
        pixel_data[18][138] = 4'b0111; // x=138, y=18
        pixel_data[18][139] = 4'b0111; // x=139, y=18
        pixel_data[18][140] = 4'b0111; // x=140, y=18
        pixel_data[18][141] = 4'b0111; // x=141, y=18
        pixel_data[18][142] = 4'b0111; // x=142, y=18
        pixel_data[18][143] = 4'b0111; // x=143, y=18
        pixel_data[18][144] = 4'b0111; // x=144, y=18
        pixel_data[18][145] = 4'b0111; // x=145, y=18
        pixel_data[18][146] = 4'b0111; // x=146, y=18
        pixel_data[18][147] = 4'b0111; // x=147, y=18
        pixel_data[18][148] = 4'b0111; // x=148, y=18
        pixel_data[18][149] = 4'b0111; // x=149, y=18
        pixel_data[18][150] = 4'b0111; // x=150, y=18
        pixel_data[18][151] = 4'b0111; // x=151, y=18
        pixel_data[18][152] = 4'b0111; // x=152, y=18
        pixel_data[18][153] = 4'b0111; // x=153, y=18
        pixel_data[18][154] = 4'b0111; // x=154, y=18
        pixel_data[18][155] = 4'b0111; // x=155, y=18
        pixel_data[18][156] = 4'b0111; // x=156, y=18
        pixel_data[18][157] = 4'b0111; // x=157, y=18
        pixel_data[18][158] = 4'b0111; // x=158, y=18
        pixel_data[18][159] = 4'b0111; // x=159, y=18
        pixel_data[18][160] = 4'b0111; // x=160, y=18
        pixel_data[18][161] = 4'b0111; // x=161, y=18
        pixel_data[18][162] = 4'b0111; // x=162, y=18
        pixel_data[18][163] = 4'b0111; // x=163, y=18
        pixel_data[18][164] = 4'b0111; // x=164, y=18
        pixel_data[18][165] = 4'b0111; // x=165, y=18
        pixel_data[18][166] = 4'b0111; // x=166, y=18
        pixel_data[18][167] = 4'b0111; // x=167, y=18
        pixel_data[18][168] = 4'b0111; // x=168, y=18
        pixel_data[18][169] = 4'b0111; // x=169, y=18
        pixel_data[18][170] = 4'b0111; // x=170, y=18
        pixel_data[18][171] = 4'b0111; // x=171, y=18
        pixel_data[18][172] = 4'b0111; // x=172, y=18
        pixel_data[18][173] = 4'b0111; // x=173, y=18
        pixel_data[18][174] = 4'b0111; // x=174, y=18
        pixel_data[18][175] = 4'b0111; // x=175, y=18
        pixel_data[18][176] = 4'b0111; // x=176, y=18
        pixel_data[18][177] = 4'b0111; // x=177, y=18
        pixel_data[18][178] = 4'b0111; // x=178, y=18
        pixel_data[18][179] = 4'b0111; // x=179, y=18
        pixel_data[19][0] = 4'b0111; // x=0, y=19
        pixel_data[19][1] = 4'b0111; // x=1, y=19
        pixel_data[19][2] = 4'b0111; // x=2, y=19
        pixel_data[19][3] = 4'b0111; // x=3, y=19
        pixel_data[19][4] = 4'b0111; // x=4, y=19
        pixel_data[19][5] = 4'b0111; // x=5, y=19
        pixel_data[19][6] = 4'b0111; // x=6, y=19
        pixel_data[19][7] = 4'b0111; // x=7, y=19
        pixel_data[19][8] = 4'b0111; // x=8, y=19
        pixel_data[19][9] = 4'b0111; // x=9, y=19
        pixel_data[19][10] = 4'b0000; // x=10, y=19
        pixel_data[19][11] = 4'b0111; // x=11, y=19
        pixel_data[19][12] = 4'b1010; // x=12, y=19
        pixel_data[19][13] = 4'b1011; // x=13, y=19
        pixel_data[19][14] = 4'b1101; // x=14, y=19
        pixel_data[19][15] = 4'b1101; // x=15, y=19
        pixel_data[19][16] = 4'b0001; // x=16, y=19
        pixel_data[19][17] = 4'b0001; // x=17, y=19
        pixel_data[19][18] = 4'b0001; // x=18, y=19
        pixel_data[19][19] = 4'b0001; // x=19, y=19
        pixel_data[19][20] = 4'b1101; // x=20, y=19
        pixel_data[19][21] = 4'b1101; // x=21, y=19
        pixel_data[19][22] = 4'b0001; // x=22, y=19
        pixel_data[19][23] = 4'b0001; // x=23, y=19
        pixel_data[19][24] = 4'b0001; // x=24, y=19
        pixel_data[19][25] = 4'b0001; // x=25, y=19
        pixel_data[19][26] = 4'b1101; // x=26, y=19
        pixel_data[19][27] = 4'b1101; // x=27, y=19
        pixel_data[19][28] = 4'b1101; // x=28, y=19
        pixel_data[19][29] = 4'b0101; // x=29, y=19
        pixel_data[19][30] = 4'b0000; // x=30, y=19
        pixel_data[19][31] = 4'b0111; // x=31, y=19
        pixel_data[19][32] = 4'b0111; // x=32, y=19
        pixel_data[19][33] = 4'b0111; // x=33, y=19
        pixel_data[19][34] = 4'b0111; // x=34, y=19
        pixel_data[19][35] = 4'b0111; // x=35, y=19
        pixel_data[19][36] = 4'b0111; // x=36, y=19
        pixel_data[19][37] = 4'b0111; // x=37, y=19
        pixel_data[19][38] = 4'b0111; // x=38, y=19
        pixel_data[19][39] = 4'b0111; // x=39, y=19
        pixel_data[19][40] = 4'b0111; // x=40, y=19
        pixel_data[19][41] = 4'b0111; // x=41, y=19
        pixel_data[19][42] = 4'b0111; // x=42, y=19
        pixel_data[19][43] = 4'b0111; // x=43, y=19
        pixel_data[19][44] = 4'b0111; // x=44, y=19
        pixel_data[19][45] = 4'b0111; // x=45, y=19
        pixel_data[19][46] = 4'b0111; // x=46, y=19
        pixel_data[19][47] = 4'b0111; // x=47, y=19
        pixel_data[19][48] = 4'b0111; // x=48, y=19
        pixel_data[19][49] = 4'b0111; // x=49, y=19
        pixel_data[19][50] = 4'b0111; // x=50, y=19
        pixel_data[19][51] = 4'b0111; // x=51, y=19
        pixel_data[19][52] = 4'b0111; // x=52, y=19
        pixel_data[19][53] = 4'b0111; // x=53, y=19
        pixel_data[19][54] = 4'b0111; // x=54, y=19
        pixel_data[19][55] = 4'b0111; // x=55, y=19
        pixel_data[19][56] = 4'b0111; // x=56, y=19
        pixel_data[19][57] = 4'b0111; // x=57, y=19
        pixel_data[19][58] = 4'b0111; // x=58, y=19
        pixel_data[19][59] = 4'b0111; // x=59, y=19
        pixel_data[19][60] = 4'b0111; // x=60, y=19
        pixel_data[19][61] = 4'b0111; // x=61, y=19
        pixel_data[19][62] = 4'b0111; // x=62, y=19
        pixel_data[19][63] = 4'b0111; // x=63, y=19
        pixel_data[19][64] = 4'b0111; // x=64, y=19
        pixel_data[19][65] = 4'b0111; // x=65, y=19
        pixel_data[19][66] = 4'b0111; // x=66, y=19
        pixel_data[19][67] = 4'b0111; // x=67, y=19
        pixel_data[19][68] = 4'b0111; // x=68, y=19
        pixel_data[19][69] = 4'b0111; // x=69, y=19
        pixel_data[19][70] = 4'b0111; // x=70, y=19
        pixel_data[19][71] = 4'b0111; // x=71, y=19
        pixel_data[19][72] = 4'b0111; // x=72, y=19
        pixel_data[19][73] = 4'b0111; // x=73, y=19
        pixel_data[19][74] = 4'b0111; // x=74, y=19
        pixel_data[19][75] = 4'b0111; // x=75, y=19
        pixel_data[19][76] = 4'b0111; // x=76, y=19
        pixel_data[19][77] = 4'b0111; // x=77, y=19
        pixel_data[19][78] = 4'b0111; // x=78, y=19
        pixel_data[19][79] = 4'b0111; // x=79, y=19
        pixel_data[19][80] = 4'b0111; // x=80, y=19
        pixel_data[19][81] = 4'b0111; // x=81, y=19
        pixel_data[19][82] = 4'b0111; // x=82, y=19
        pixel_data[19][83] = 4'b0111; // x=83, y=19
        pixel_data[19][84] = 4'b0111; // x=84, y=19
        pixel_data[19][85] = 4'b0111; // x=85, y=19
        pixel_data[19][86] = 4'b0111; // x=86, y=19
        pixel_data[19][87] = 4'b0111; // x=87, y=19
        pixel_data[19][88] = 4'b0111; // x=88, y=19
        pixel_data[19][89] = 4'b0111; // x=89, y=19
        pixel_data[19][90] = 4'b0111; // x=90, y=19
        pixel_data[19][91] = 4'b0111; // x=91, y=19
        pixel_data[19][92] = 4'b0111; // x=92, y=19
        pixel_data[19][93] = 4'b0111; // x=93, y=19
        pixel_data[19][94] = 4'b0111; // x=94, y=19
        pixel_data[19][95] = 4'b0111; // x=95, y=19
        pixel_data[19][96] = 4'b0111; // x=96, y=19
        pixel_data[19][97] = 4'b0111; // x=97, y=19
        pixel_data[19][98] = 4'b0111; // x=98, y=19
        pixel_data[19][99] = 4'b0111; // x=99, y=19
        pixel_data[19][100] = 4'b0111; // x=100, y=19
        pixel_data[19][101] = 4'b0111; // x=101, y=19
        pixel_data[19][102] = 4'b0111; // x=102, y=19
        pixel_data[19][103] = 4'b0111; // x=103, y=19
        pixel_data[19][104] = 4'b0111; // x=104, y=19
        pixel_data[19][105] = 4'b0111; // x=105, y=19
        pixel_data[19][106] = 4'b0111; // x=106, y=19
        pixel_data[19][107] = 4'b0111; // x=107, y=19
        pixel_data[19][108] = 4'b0111; // x=108, y=19
        pixel_data[19][109] = 4'b0111; // x=109, y=19
        pixel_data[19][110] = 4'b0111; // x=110, y=19
        pixel_data[19][111] = 4'b0111; // x=111, y=19
        pixel_data[19][112] = 4'b0111; // x=112, y=19
        pixel_data[19][113] = 4'b0111; // x=113, y=19
        pixel_data[19][114] = 4'b0111; // x=114, y=19
        pixel_data[19][115] = 4'b0111; // x=115, y=19
        pixel_data[19][116] = 4'b0111; // x=116, y=19
        pixel_data[19][117] = 4'b0111; // x=117, y=19
        pixel_data[19][118] = 4'b0111; // x=118, y=19
        pixel_data[19][119] = 4'b0111; // x=119, y=19
        pixel_data[19][120] = 4'b0111; // x=120, y=19
        pixel_data[19][121] = 4'b0111; // x=121, y=19
        pixel_data[19][122] = 4'b0111; // x=122, y=19
        pixel_data[19][123] = 4'b0111; // x=123, y=19
        pixel_data[19][124] = 4'b0111; // x=124, y=19
        pixel_data[19][125] = 4'b0111; // x=125, y=19
        pixel_data[19][126] = 4'b0111; // x=126, y=19
        pixel_data[19][127] = 4'b0111; // x=127, y=19
        pixel_data[19][128] = 4'b0111; // x=128, y=19
        pixel_data[19][129] = 4'b0111; // x=129, y=19
        pixel_data[19][130] = 4'b0111; // x=130, y=19
        pixel_data[19][131] = 4'b0111; // x=131, y=19
        pixel_data[19][132] = 4'b0111; // x=132, y=19
        pixel_data[19][133] = 4'b0111; // x=133, y=19
        pixel_data[19][134] = 4'b0111; // x=134, y=19
        pixel_data[19][135] = 4'b0111; // x=135, y=19
        pixel_data[19][136] = 4'b0111; // x=136, y=19
        pixel_data[19][137] = 4'b0111; // x=137, y=19
        pixel_data[19][138] = 4'b0111; // x=138, y=19
        pixel_data[19][139] = 4'b0111; // x=139, y=19
        pixel_data[19][140] = 4'b0111; // x=140, y=19
        pixel_data[19][141] = 4'b0111; // x=141, y=19
        pixel_data[19][142] = 4'b0111; // x=142, y=19
        pixel_data[19][143] = 4'b0111; // x=143, y=19
        pixel_data[19][144] = 4'b0111; // x=144, y=19
        pixel_data[19][145] = 4'b0111; // x=145, y=19
        pixel_data[19][146] = 4'b0111; // x=146, y=19
        pixel_data[19][147] = 4'b0111; // x=147, y=19
        pixel_data[19][148] = 4'b0111; // x=148, y=19
        pixel_data[19][149] = 4'b0111; // x=149, y=19
        pixel_data[19][150] = 4'b0111; // x=150, y=19
        pixel_data[19][151] = 4'b0111; // x=151, y=19
        pixel_data[19][152] = 4'b0111; // x=152, y=19
        pixel_data[19][153] = 4'b0111; // x=153, y=19
        pixel_data[19][154] = 4'b0111; // x=154, y=19
        pixel_data[19][155] = 4'b0111; // x=155, y=19
        pixel_data[19][156] = 4'b0111; // x=156, y=19
        pixel_data[19][157] = 4'b0111; // x=157, y=19
        pixel_data[19][158] = 4'b0111; // x=158, y=19
        pixel_data[19][159] = 4'b0111; // x=159, y=19
        pixel_data[19][160] = 4'b0111; // x=160, y=19
        pixel_data[19][161] = 4'b0111; // x=161, y=19
        pixel_data[19][162] = 4'b0111; // x=162, y=19
        pixel_data[19][163] = 4'b0111; // x=163, y=19
        pixel_data[19][164] = 4'b0111; // x=164, y=19
        pixel_data[19][165] = 4'b0111; // x=165, y=19
        pixel_data[19][166] = 4'b0111; // x=166, y=19
        pixel_data[19][167] = 4'b0111; // x=167, y=19
        pixel_data[19][168] = 4'b0111; // x=168, y=19
        pixel_data[19][169] = 4'b0111; // x=169, y=19
        pixel_data[19][170] = 4'b0111; // x=170, y=19
        pixel_data[19][171] = 4'b0111; // x=171, y=19
        pixel_data[19][172] = 4'b0111; // x=172, y=19
        pixel_data[19][173] = 4'b0111; // x=173, y=19
        pixel_data[19][174] = 4'b0111; // x=174, y=19
        pixel_data[19][175] = 4'b0111; // x=175, y=19
        pixel_data[19][176] = 4'b0111; // x=176, y=19
        pixel_data[19][177] = 4'b0111; // x=177, y=19
        pixel_data[19][178] = 4'b0111; // x=178, y=19
        pixel_data[19][179] = 4'b0111; // x=179, y=19
        pixel_data[20][0] = 4'b0111; // x=0, y=20
        pixel_data[20][1] = 4'b0111; // x=1, y=20
        pixel_data[20][2] = 4'b0111; // x=2, y=20
        pixel_data[20][3] = 4'b0111; // x=3, y=20
        pixel_data[20][4] = 4'b0111; // x=4, y=20
        pixel_data[20][5] = 4'b0111; // x=5, y=20
        pixel_data[20][6] = 4'b0111; // x=6, y=20
        pixel_data[20][7] = 4'b0111; // x=7, y=20
        pixel_data[20][8] = 4'b0111; // x=8, y=20
        pixel_data[20][9] = 4'b0000; // x=9, y=20
        pixel_data[20][10] = 4'b0111; // x=10, y=20
        pixel_data[20][11] = 4'b0010; // x=11, y=20
        pixel_data[20][12] = 4'b1101; // x=12, y=20
        pixel_data[20][13] = 4'b1101; // x=13, y=20
        pixel_data[20][14] = 4'b0001; // x=14, y=20
        pixel_data[20][15] = 4'b0001; // x=15, y=20
        pixel_data[20][16] = 4'b0001; // x=16, y=20
        pixel_data[20][17] = 4'b1101; // x=17, y=20
        pixel_data[20][18] = 4'b1101; // x=18, y=20
        pixel_data[20][19] = 4'b1101; // x=19, y=20
        pixel_data[20][20] = 4'b0001; // x=20, y=20
        pixel_data[20][21] = 4'b0001; // x=21, y=20
        pixel_data[20][22] = 4'b1101; // x=22, y=20
        pixel_data[20][23] = 4'b1101; // x=23, y=20
        pixel_data[20][24] = 4'b1101; // x=24, y=20
        pixel_data[20][25] = 4'b0001; // x=25, y=20
        pixel_data[20][26] = 4'b0001; // x=26, y=20
        pixel_data[20][27] = 4'b0001; // x=27, y=20
        pixel_data[20][28] = 4'b0001; // x=28, y=20
        pixel_data[20][29] = 4'b1101; // x=29, y=20
        pixel_data[20][30] = 4'b1100; // x=30, y=20
        pixel_data[20][31] = 4'b1110; // x=31, y=20
        pixel_data[20][32] = 4'b0111; // x=32, y=20
        pixel_data[20][33] = 4'b0111; // x=33, y=20
        pixel_data[20][34] = 4'b0111; // x=34, y=20
        pixel_data[20][35] = 4'b0111; // x=35, y=20
        pixel_data[20][36] = 4'b0111; // x=36, y=20
        pixel_data[20][37] = 4'b0111; // x=37, y=20
        pixel_data[20][38] = 4'b0111; // x=38, y=20
        pixel_data[20][39] = 4'b0111; // x=39, y=20
        pixel_data[20][40] = 4'b0111; // x=40, y=20
        pixel_data[20][41] = 4'b0111; // x=41, y=20
        pixel_data[20][42] = 4'b0111; // x=42, y=20
        pixel_data[20][43] = 4'b0111; // x=43, y=20
        pixel_data[20][44] = 4'b0111; // x=44, y=20
        pixel_data[20][45] = 4'b0111; // x=45, y=20
        pixel_data[20][46] = 4'b0111; // x=46, y=20
        pixel_data[20][47] = 4'b0111; // x=47, y=20
        pixel_data[20][48] = 4'b0111; // x=48, y=20
        pixel_data[20][49] = 4'b0111; // x=49, y=20
        pixel_data[20][50] = 4'b0111; // x=50, y=20
        pixel_data[20][51] = 4'b0111; // x=51, y=20
        pixel_data[20][52] = 4'b0111; // x=52, y=20
        pixel_data[20][53] = 4'b0111; // x=53, y=20
        pixel_data[20][54] = 4'b0111; // x=54, y=20
        pixel_data[20][55] = 4'b0111; // x=55, y=20
        pixel_data[20][56] = 4'b0111; // x=56, y=20
        pixel_data[20][57] = 4'b0111; // x=57, y=20
        pixel_data[20][58] = 4'b0111; // x=58, y=20
        pixel_data[20][59] = 4'b0111; // x=59, y=20
        pixel_data[20][60] = 4'b0111; // x=60, y=20
        pixel_data[20][61] = 4'b0111; // x=61, y=20
        pixel_data[20][62] = 4'b0111; // x=62, y=20
        pixel_data[20][63] = 4'b0111; // x=63, y=20
        pixel_data[20][64] = 4'b0111; // x=64, y=20
        pixel_data[20][65] = 4'b0111; // x=65, y=20
        pixel_data[20][66] = 4'b0111; // x=66, y=20
        pixel_data[20][67] = 4'b0111; // x=67, y=20
        pixel_data[20][68] = 4'b0111; // x=68, y=20
        pixel_data[20][69] = 4'b0111; // x=69, y=20
        pixel_data[20][70] = 4'b0111; // x=70, y=20
        pixel_data[20][71] = 4'b0111; // x=71, y=20
        pixel_data[20][72] = 4'b0111; // x=72, y=20
        pixel_data[20][73] = 4'b0111; // x=73, y=20
        pixel_data[20][74] = 4'b0111; // x=74, y=20
        pixel_data[20][75] = 4'b0111; // x=75, y=20
        pixel_data[20][76] = 4'b0111; // x=76, y=20
        pixel_data[20][77] = 4'b0111; // x=77, y=20
        pixel_data[20][78] = 4'b0111; // x=78, y=20
        pixel_data[20][79] = 4'b0111; // x=79, y=20
        pixel_data[20][80] = 4'b0111; // x=80, y=20
        pixel_data[20][81] = 4'b0111; // x=81, y=20
        pixel_data[20][82] = 4'b0111; // x=82, y=20
        pixel_data[20][83] = 4'b0111; // x=83, y=20
        pixel_data[20][84] = 4'b0111; // x=84, y=20
        pixel_data[20][85] = 4'b0111; // x=85, y=20
        pixel_data[20][86] = 4'b0111; // x=86, y=20
        pixel_data[20][87] = 4'b0111; // x=87, y=20
        pixel_data[20][88] = 4'b0111; // x=88, y=20
        pixel_data[20][89] = 4'b0111; // x=89, y=20
        pixel_data[20][90] = 4'b0111; // x=90, y=20
        pixel_data[20][91] = 4'b0111; // x=91, y=20
        pixel_data[20][92] = 4'b0111; // x=92, y=20
        pixel_data[20][93] = 4'b0111; // x=93, y=20
        pixel_data[20][94] = 4'b0111; // x=94, y=20
        pixel_data[20][95] = 4'b0111; // x=95, y=20
        pixel_data[20][96] = 4'b0111; // x=96, y=20
        pixel_data[20][97] = 4'b0111; // x=97, y=20
        pixel_data[20][98] = 4'b0111; // x=98, y=20
        pixel_data[20][99] = 4'b0111; // x=99, y=20
        pixel_data[20][100] = 4'b0111; // x=100, y=20
        pixel_data[20][101] = 4'b0111; // x=101, y=20
        pixel_data[20][102] = 4'b0111; // x=102, y=20
        pixel_data[20][103] = 4'b0111; // x=103, y=20
        pixel_data[20][104] = 4'b0111; // x=104, y=20
        pixel_data[20][105] = 4'b0111; // x=105, y=20
        pixel_data[20][106] = 4'b0111; // x=106, y=20
        pixel_data[20][107] = 4'b0111; // x=107, y=20
        pixel_data[20][108] = 4'b0111; // x=108, y=20
        pixel_data[20][109] = 4'b0111; // x=109, y=20
        pixel_data[20][110] = 4'b0111; // x=110, y=20
        pixel_data[20][111] = 4'b0111; // x=111, y=20
        pixel_data[20][112] = 4'b0111; // x=112, y=20
        pixel_data[20][113] = 4'b0111; // x=113, y=20
        pixel_data[20][114] = 4'b0111; // x=114, y=20
        pixel_data[20][115] = 4'b0111; // x=115, y=20
        pixel_data[20][116] = 4'b0111; // x=116, y=20
        pixel_data[20][117] = 4'b0111; // x=117, y=20
        pixel_data[20][118] = 4'b0111; // x=118, y=20
        pixel_data[20][119] = 4'b0111; // x=119, y=20
        pixel_data[20][120] = 4'b0111; // x=120, y=20
        pixel_data[20][121] = 4'b0111; // x=121, y=20
        pixel_data[20][122] = 4'b0111; // x=122, y=20
        pixel_data[20][123] = 4'b0111; // x=123, y=20
        pixel_data[20][124] = 4'b0111; // x=124, y=20
        pixel_data[20][125] = 4'b0111; // x=125, y=20
        pixel_data[20][126] = 4'b0111; // x=126, y=20
        pixel_data[20][127] = 4'b0111; // x=127, y=20
        pixel_data[20][128] = 4'b0111; // x=128, y=20
        pixel_data[20][129] = 4'b0111; // x=129, y=20
        pixel_data[20][130] = 4'b0111; // x=130, y=20
        pixel_data[20][131] = 4'b0111; // x=131, y=20
        pixel_data[20][132] = 4'b0111; // x=132, y=20
        pixel_data[20][133] = 4'b0111; // x=133, y=20
        pixel_data[20][134] = 4'b0111; // x=134, y=20
        pixel_data[20][135] = 4'b0111; // x=135, y=20
        pixel_data[20][136] = 4'b0111; // x=136, y=20
        pixel_data[20][137] = 4'b0111; // x=137, y=20
        pixel_data[20][138] = 4'b0111; // x=138, y=20
        pixel_data[20][139] = 4'b0111; // x=139, y=20
        pixel_data[20][140] = 4'b0111; // x=140, y=20
        pixel_data[20][141] = 4'b0111; // x=141, y=20
        pixel_data[20][142] = 4'b0111; // x=142, y=20
        pixel_data[20][143] = 4'b0111; // x=143, y=20
        pixel_data[20][144] = 4'b0111; // x=144, y=20
        pixel_data[20][145] = 4'b0111; // x=145, y=20
        pixel_data[20][146] = 4'b0111; // x=146, y=20
        pixel_data[20][147] = 4'b0111; // x=147, y=20
        pixel_data[20][148] = 4'b0111; // x=148, y=20
        pixel_data[20][149] = 4'b0111; // x=149, y=20
        pixel_data[20][150] = 4'b0111; // x=150, y=20
        pixel_data[20][151] = 4'b0111; // x=151, y=20
        pixel_data[20][152] = 4'b0111; // x=152, y=20
        pixel_data[20][153] = 4'b0111; // x=153, y=20
        pixel_data[20][154] = 4'b0111; // x=154, y=20
        pixel_data[20][155] = 4'b0111; // x=155, y=20
        pixel_data[20][156] = 4'b0111; // x=156, y=20
        pixel_data[20][157] = 4'b0111; // x=157, y=20
        pixel_data[20][158] = 4'b0111; // x=158, y=20
        pixel_data[20][159] = 4'b0111; // x=159, y=20
        pixel_data[20][160] = 4'b0111; // x=160, y=20
        pixel_data[20][161] = 4'b0111; // x=161, y=20
        pixel_data[20][162] = 4'b0111; // x=162, y=20
        pixel_data[20][163] = 4'b0111; // x=163, y=20
        pixel_data[20][164] = 4'b0111; // x=164, y=20
        pixel_data[20][165] = 4'b0111; // x=165, y=20
        pixel_data[20][166] = 4'b0111; // x=166, y=20
        pixel_data[20][167] = 4'b0111; // x=167, y=20
        pixel_data[20][168] = 4'b0111; // x=168, y=20
        pixel_data[20][169] = 4'b0111; // x=169, y=20
        pixel_data[20][170] = 4'b0111; // x=170, y=20
        pixel_data[20][171] = 4'b0111; // x=171, y=20
        pixel_data[20][172] = 4'b0111; // x=172, y=20
        pixel_data[20][173] = 4'b0111; // x=173, y=20
        pixel_data[20][174] = 4'b0111; // x=174, y=20
        pixel_data[20][175] = 4'b0111; // x=175, y=20
        pixel_data[20][176] = 4'b0111; // x=176, y=20
        pixel_data[20][177] = 4'b0111; // x=177, y=20
        pixel_data[20][178] = 4'b0111; // x=178, y=20
        pixel_data[20][179] = 4'b0111; // x=179, y=20
        pixel_data[21][0] = 4'b0111; // x=0, y=21
        pixel_data[21][1] = 4'b0111; // x=1, y=21
        pixel_data[21][2] = 4'b0111; // x=2, y=21
        pixel_data[21][3] = 4'b0111; // x=3, y=21
        pixel_data[21][4] = 4'b0111; // x=4, y=21
        pixel_data[21][5] = 4'b0111; // x=5, y=21
        pixel_data[21][6] = 4'b0111; // x=6, y=21
        pixel_data[21][7] = 4'b0111; // x=7, y=21
        pixel_data[21][8] = 4'b0111; // x=8, y=21
        pixel_data[21][9] = 4'b0111; // x=9, y=21
        pixel_data[21][10] = 4'b0100; // x=10, y=21
        pixel_data[21][11] = 4'b1101; // x=11, y=21
        pixel_data[21][12] = 4'b1101; // x=12, y=21
        pixel_data[21][13] = 4'b1101; // x=13, y=21
        pixel_data[21][14] = 4'b0001; // x=14, y=21
        pixel_data[21][15] = 4'b1101; // x=15, y=21
        pixel_data[21][16] = 4'b1101; // x=16, y=21
        pixel_data[21][17] = 4'b1111; // x=17, y=21
        pixel_data[21][18] = 4'b1001; // x=18, y=21
        pixel_data[21][19] = 4'b0100; // x=19, y=21
        pixel_data[21][20] = 4'b0110; // x=20, y=21
        pixel_data[21][21] = 4'b0110; // x=21, y=21
        pixel_data[21][22] = 4'b0100; // x=22, y=21
        pixel_data[21][23] = 4'b0010; // x=23, y=21
        pixel_data[21][24] = 4'b0011; // x=24, y=21
        pixel_data[21][25] = 4'b1101; // x=25, y=21
        pixel_data[21][26] = 4'b1101; // x=26, y=21
        pixel_data[21][27] = 4'b0001; // x=27, y=21
        pixel_data[21][28] = 4'b0001; // x=28, y=21
        pixel_data[21][29] = 4'b1101; // x=29, y=21
        pixel_data[21][30] = 4'b1101; // x=30, y=21
        pixel_data[21][31] = 4'b0100; // x=31, y=21
        pixel_data[21][32] = 4'b0111; // x=32, y=21
        pixel_data[21][33] = 4'b0000; // x=33, y=21
        pixel_data[21][34] = 4'b0111; // x=34, y=21
        pixel_data[21][35] = 4'b0111; // x=35, y=21
        pixel_data[21][36] = 4'b0111; // x=36, y=21
        pixel_data[21][37] = 4'b0111; // x=37, y=21
        pixel_data[21][38] = 4'b0111; // x=38, y=21
        pixel_data[21][39] = 4'b0111; // x=39, y=21
        pixel_data[21][40] = 4'b0111; // x=40, y=21
        pixel_data[21][41] = 4'b0111; // x=41, y=21
        pixel_data[21][42] = 4'b0000; // x=42, y=21
        pixel_data[21][43] = 4'b0000; // x=43, y=21
        pixel_data[21][44] = 4'b0000; // x=44, y=21
        pixel_data[21][45] = 4'b0000; // x=45, y=21
        pixel_data[21][46] = 4'b0111; // x=46, y=21
        pixel_data[21][47] = 4'b0111; // x=47, y=21
        pixel_data[21][48] = 4'b0111; // x=48, y=21
        pixel_data[21][49] = 4'b0000; // x=49, y=21
        pixel_data[21][50] = 4'b0000; // x=50, y=21
        pixel_data[21][51] = 4'b0000; // x=51, y=21
        pixel_data[21][52] = 4'b0000; // x=52, y=21
        pixel_data[21][53] = 4'b0000; // x=53, y=21
        pixel_data[21][54] = 4'b0111; // x=54, y=21
        pixel_data[21][55] = 4'b0111; // x=55, y=21
        pixel_data[21][56] = 4'b0111; // x=56, y=21
        pixel_data[21][57] = 4'b0111; // x=57, y=21
        pixel_data[21][58] = 4'b0111; // x=58, y=21
        pixel_data[21][59] = 4'b0111; // x=59, y=21
        pixel_data[21][60] = 4'b0111; // x=60, y=21
        pixel_data[21][61] = 4'b0111; // x=61, y=21
        pixel_data[21][62] = 4'b0111; // x=62, y=21
        pixel_data[21][63] = 4'b0111; // x=63, y=21
        pixel_data[21][64] = 4'b0111; // x=64, y=21
        pixel_data[21][65] = 4'b0000; // x=65, y=21
        pixel_data[21][66] = 4'b0000; // x=66, y=21
        pixel_data[21][67] = 4'b0000; // x=67, y=21
        pixel_data[21][68] = 4'b0000; // x=68, y=21
        pixel_data[21][69] = 4'b0111; // x=69, y=21
        pixel_data[21][70] = 4'b0111; // x=70, y=21
        pixel_data[21][71] = 4'b0111; // x=71, y=21
        pixel_data[21][72] = 4'b0000; // x=72, y=21
        pixel_data[21][73] = 4'b0000; // x=73, y=21
        pixel_data[21][74] = 4'b0000; // x=74, y=21
        pixel_data[21][75] = 4'b0000; // x=75, y=21
        pixel_data[21][76] = 4'b0111; // x=76, y=21
        pixel_data[21][77] = 4'b0111; // x=77, y=21
        pixel_data[21][78] = 4'b0111; // x=78, y=21
        pixel_data[21][79] = 4'b0111; // x=79, y=21
        pixel_data[21][80] = 4'b0111; // x=80, y=21
        pixel_data[21][81] = 4'b0111; // x=81, y=21
        pixel_data[21][82] = 4'b0111; // x=82, y=21
        pixel_data[21][83] = 4'b0111; // x=83, y=21
        pixel_data[21][84] = 4'b0111; // x=84, y=21
        pixel_data[21][85] = 4'b0111; // x=85, y=21
        pixel_data[21][86] = 4'b0111; // x=86, y=21
        pixel_data[21][87] = 4'b0000; // x=87, y=21
        pixel_data[21][88] = 4'b0000; // x=88, y=21
        pixel_data[21][89] = 4'b0000; // x=89, y=21
        pixel_data[21][90] = 4'b0000; // x=90, y=21
        pixel_data[21][91] = 4'b0000; // x=91, y=21
        pixel_data[21][92] = 4'b0000; // x=92, y=21
        pixel_data[21][93] = 4'b0111; // x=93, y=21
        pixel_data[21][94] = 4'b0111; // x=94, y=21
        pixel_data[21][95] = 4'b0111; // x=95, y=21
        pixel_data[21][96] = 4'b0000; // x=96, y=21
        pixel_data[21][97] = 4'b0000; // x=97, y=21
        pixel_data[21][98] = 4'b0000; // x=98, y=21
        pixel_data[21][99] = 4'b0000; // x=99, y=21
        pixel_data[21][100] = 4'b0111; // x=100, y=21
        pixel_data[21][101] = 4'b0111; // x=101, y=21
        pixel_data[21][102] = 4'b0000; // x=102, y=21
        pixel_data[21][103] = 4'b0111; // x=103, y=21
        pixel_data[21][104] = 4'b0111; // x=104, y=21
        pixel_data[21][105] = 4'b0111; // x=105, y=21
        pixel_data[21][106] = 4'b0111; // x=106, y=21
        pixel_data[21][107] = 4'b0111; // x=107, y=21
        pixel_data[21][108] = 4'b0111; // x=108, y=21
        pixel_data[21][109] = 4'b0111; // x=109, y=21
        pixel_data[21][110] = 4'b0000; // x=110, y=21
        pixel_data[21][111] = 4'b0000; // x=111, y=21
        pixel_data[21][112] = 4'b0000; // x=112, y=21
        pixel_data[21][113] = 4'b0111; // x=113, y=21
        pixel_data[21][114] = 4'b0111; // x=114, y=21
        pixel_data[21][115] = 4'b0111; // x=115, y=21
        pixel_data[21][116] = 4'b0111; // x=116, y=21
        pixel_data[21][117] = 4'b0111; // x=117, y=21
        pixel_data[21][118] = 4'b0000; // x=118, y=21
        pixel_data[21][119] = 4'b0000; // x=119, y=21
        pixel_data[21][120] = 4'b0000; // x=120, y=21
        pixel_data[21][121] = 4'b0111; // x=121, y=21
        pixel_data[21][122] = 4'b0111; // x=122, y=21
        pixel_data[21][123] = 4'b0111; // x=123, y=21
        pixel_data[21][124] = 4'b0111; // x=124, y=21
        pixel_data[21][125] = 4'b0111; // x=125, y=21
        pixel_data[21][126] = 4'b0111; // x=126, y=21
        pixel_data[21][127] = 4'b0111; // x=127, y=21
        pixel_data[21][128] = 4'b0111; // x=128, y=21
        pixel_data[21][129] = 4'b0111; // x=129, y=21
        pixel_data[21][130] = 4'b0111; // x=130, y=21
        pixel_data[21][131] = 4'b0111; // x=131, y=21
        pixel_data[21][132] = 4'b0111; // x=132, y=21
        pixel_data[21][133] = 4'b0111; // x=133, y=21
        pixel_data[21][134] = 4'b0111; // x=134, y=21
        pixel_data[21][135] = 4'b0111; // x=135, y=21
        pixel_data[21][136] = 4'b0111; // x=136, y=21
        pixel_data[21][137] = 4'b0111; // x=137, y=21
        pixel_data[21][138] = 4'b0111; // x=138, y=21
        pixel_data[21][139] = 4'b0111; // x=139, y=21
        pixel_data[21][140] = 4'b0111; // x=140, y=21
        pixel_data[21][141] = 4'b0111; // x=141, y=21
        pixel_data[21][142] = 4'b0111; // x=142, y=21
        pixel_data[21][143] = 4'b0000; // x=143, y=21
        pixel_data[21][144] = 4'b0000; // x=144, y=21
        pixel_data[21][145] = 4'b0111; // x=145, y=21
        pixel_data[21][146] = 4'b0111; // x=146, y=21
        pixel_data[21][147] = 4'b0000; // x=147, y=21
        pixel_data[21][148] = 4'b0000; // x=148, y=21
        pixel_data[21][149] = 4'b0111; // x=149, y=21
        pixel_data[21][150] = 4'b0111; // x=150, y=21
        pixel_data[21][151] = 4'b0111; // x=151, y=21
        pixel_data[21][152] = 4'b0111; // x=152, y=21
        pixel_data[21][153] = 4'b0111; // x=153, y=21
        pixel_data[21][154] = 4'b0111; // x=154, y=21
        pixel_data[21][155] = 4'b0111; // x=155, y=21
        pixel_data[21][156] = 4'b0111; // x=156, y=21
        pixel_data[21][157] = 4'b0111; // x=157, y=21
        pixel_data[21][158] = 4'b0111; // x=158, y=21
        pixel_data[21][159] = 4'b0111; // x=159, y=21
        pixel_data[21][160] = 4'b0111; // x=160, y=21
        pixel_data[21][161] = 4'b0111; // x=161, y=21
        pixel_data[21][162] = 4'b0111; // x=162, y=21
        pixel_data[21][163] = 4'b0111; // x=163, y=21
        pixel_data[21][164] = 4'b0111; // x=164, y=21
        pixel_data[21][165] = 4'b0111; // x=165, y=21
        pixel_data[21][166] = 4'b0111; // x=166, y=21
        pixel_data[21][167] = 4'b0111; // x=167, y=21
        pixel_data[21][168] = 4'b0111; // x=168, y=21
        pixel_data[21][169] = 4'b0111; // x=169, y=21
        pixel_data[21][170] = 4'b0111; // x=170, y=21
        pixel_data[21][171] = 4'b0111; // x=171, y=21
        pixel_data[21][172] = 4'b0111; // x=172, y=21
        pixel_data[21][173] = 4'b0111; // x=173, y=21
        pixel_data[21][174] = 4'b0111; // x=174, y=21
        pixel_data[21][175] = 4'b0111; // x=175, y=21
        pixel_data[21][176] = 4'b0111; // x=176, y=21
        pixel_data[21][177] = 4'b0111; // x=177, y=21
        pixel_data[21][178] = 4'b0111; // x=178, y=21
        pixel_data[21][179] = 4'b0111; // x=179, y=21
        pixel_data[22][0] = 4'b0111; // x=0, y=22
        pixel_data[22][1] = 4'b0111; // x=1, y=22
        pixel_data[22][2] = 4'b0111; // x=2, y=22
        pixel_data[22][3] = 4'b0111; // x=3, y=22
        pixel_data[22][4] = 4'b0111; // x=4, y=22
        pixel_data[22][5] = 4'b0111; // x=5, y=22
        pixel_data[22][6] = 4'b0111; // x=6, y=22
        pixel_data[22][7] = 4'b0111; // x=7, y=22
        pixel_data[22][8] = 4'b0111; // x=8, y=22
        pixel_data[22][9] = 4'b0111; // x=9, y=22
        pixel_data[22][10] = 4'b1000; // x=10, y=22
        pixel_data[22][11] = 4'b1101; // x=11, y=22
        pixel_data[22][12] = 4'b0001; // x=12, y=22
        pixel_data[22][13] = 4'b1101; // x=13, y=22
        pixel_data[22][14] = 4'b0001; // x=14, y=22
        pixel_data[22][15] = 4'b0001; // x=15, y=22
        pixel_data[22][16] = 4'b1001; // x=16, y=22
        pixel_data[22][17] = 4'b0111; // x=17, y=22
        pixel_data[22][18] = 4'b0111; // x=18, y=22
        pixel_data[22][19] = 4'b0111; // x=19, y=22
        pixel_data[22][20] = 4'b0111; // x=20, y=22
        pixel_data[22][21] = 4'b0111; // x=21, y=22
        pixel_data[22][22] = 4'b0111; // x=22, y=22
        pixel_data[22][23] = 4'b0111; // x=23, y=22
        pixel_data[22][24] = 4'b0000; // x=24, y=22
        pixel_data[22][25] = 4'b1001; // x=25, y=22
        pixel_data[22][26] = 4'b0011; // x=26, y=22
        pixel_data[22][27] = 4'b1101; // x=27, y=22
        pixel_data[22][28] = 4'b1101; // x=28, y=22
        pixel_data[22][29] = 4'b0011; // x=29, y=22
        pixel_data[22][30] = 4'b0100; // x=30, y=22
        pixel_data[22][31] = 4'b0111; // x=31, y=22
        pixel_data[22][32] = 4'b0111; // x=32, y=22
        pixel_data[22][33] = 4'b0111; // x=33, y=22
        pixel_data[22][34] = 4'b0111; // x=34, y=22
        pixel_data[22][35] = 4'b0111; // x=35, y=22
        pixel_data[22][36] = 4'b0111; // x=36, y=22
        pixel_data[22][37] = 4'b0111; // x=37, y=22
        pixel_data[22][38] = 4'b0111; // x=38, y=22
        pixel_data[22][39] = 4'b0111; // x=39, y=22
        pixel_data[22][40] = 4'b0000; // x=40, y=22
        pixel_data[22][41] = 4'b0000; // x=41, y=22
        pixel_data[22][42] = 4'b0111; // x=42, y=22
        pixel_data[22][43] = 4'b0111; // x=43, y=22
        pixel_data[22][44] = 4'b0111; // x=44, y=22
        pixel_data[22][45] = 4'b0111; // x=45, y=22
        pixel_data[22][46] = 4'b0111; // x=46, y=22
        pixel_data[22][47] = 4'b0000; // x=47, y=22
        pixel_data[22][48] = 4'b0111; // x=48, y=22
        pixel_data[22][49] = 4'b0111; // x=49, y=22
        pixel_data[22][50] = 4'b0111; // x=50, y=22
        pixel_data[22][51] = 4'b0111; // x=51, y=22
        pixel_data[22][52] = 4'b0111; // x=52, y=22
        pixel_data[22][53] = 4'b0000; // x=53, y=22
        pixel_data[22][54] = 4'b0000; // x=54, y=22
        pixel_data[22][55] = 4'b0111; // x=55, y=22
        pixel_data[22][56] = 4'b0111; // x=56, y=22
        pixel_data[22][57] = 4'b0111; // x=57, y=22
        pixel_data[22][58] = 4'b0111; // x=58, y=22
        pixel_data[22][59] = 4'b0111; // x=59, y=22
        pixel_data[22][60] = 4'b0111; // x=60, y=22
        pixel_data[22][61] = 4'b0111; // x=61, y=22
        pixel_data[22][62] = 4'b0111; // x=62, y=22
        pixel_data[22][63] = 4'b0000; // x=63, y=22
        pixel_data[22][64] = 4'b0000; // x=64, y=22
        pixel_data[22][65] = 4'b0000; // x=65, y=22
        pixel_data[22][66] = 4'b0111; // x=66, y=22
        pixel_data[22][67] = 4'b0111; // x=67, y=22
        pixel_data[22][68] = 4'b0111; // x=68, y=22
        pixel_data[22][69] = 4'b0111; // x=69, y=22
        pixel_data[22][70] = 4'b0000; // x=70, y=22
        pixel_data[22][71] = 4'b0000; // x=71, y=22
        pixel_data[22][72] = 4'b0111; // x=72, y=22
        pixel_data[22][73] = 4'b0111; // x=73, y=22
        pixel_data[22][74] = 4'b0111; // x=74, y=22
        pixel_data[22][75] = 4'b0111; // x=75, y=22
        pixel_data[22][76] = 4'b0111; // x=76, y=22
        pixel_data[22][77] = 4'b0000; // x=77, y=22
        pixel_data[22][78] = 4'b0000; // x=78, y=22
        pixel_data[22][79] = 4'b0111; // x=79, y=22
        pixel_data[22][80] = 4'b0111; // x=80, y=22
        pixel_data[22][81] = 4'b0111; // x=81, y=22
        pixel_data[22][82] = 4'b0111; // x=82, y=22
        pixel_data[22][83] = 4'b0111; // x=83, y=22
        pixel_data[22][84] = 4'b0111; // x=84, y=22
        pixel_data[22][85] = 4'b0000; // x=85, y=22
        pixel_data[22][86] = 4'b0000; // x=86, y=22
        pixel_data[22][87] = 4'b0111; // x=87, y=22
        pixel_data[22][88] = 4'b0111; // x=88, y=22
        pixel_data[22][89] = 4'b0111; // x=89, y=22
        pixel_data[22][90] = 4'b0111; // x=90, y=22
        pixel_data[22][91] = 4'b0111; // x=91, y=22
        pixel_data[22][92] = 4'b0111; // x=92, y=22
        pixel_data[22][93] = 4'b0111; // x=93, y=22
        pixel_data[22][94] = 4'b0000; // x=94, y=22
        pixel_data[22][95] = 4'b0000; // x=95, y=22
        pixel_data[22][96] = 4'b0111; // x=96, y=22
        pixel_data[22][97] = 4'b0111; // x=97, y=22
        pixel_data[22][98] = 4'b0111; // x=98, y=22
        pixel_data[22][99] = 4'b0000; // x=99, y=22
        pixel_data[22][100] = 4'b0000; // x=100, y=22
        pixel_data[22][101] = 4'b0111; // x=101, y=22
        pixel_data[22][102] = 4'b0111; // x=102, y=22
        pixel_data[22][103] = 4'b0111; // x=103, y=22
        pixel_data[22][104] = 4'b0111; // x=104, y=22
        pixel_data[22][105] = 4'b0111; // x=105, y=22
        pixel_data[22][106] = 4'b0111; // x=106, y=22
        pixel_data[22][107] = 4'b0111; // x=107, y=22
        pixel_data[22][108] = 4'b0000; // x=108, y=22
        pixel_data[22][109] = 4'b0111; // x=109, y=22
        pixel_data[22][110] = 4'b0111; // x=110, y=22
        pixel_data[22][111] = 4'b0111; // x=111, y=22
        pixel_data[22][112] = 4'b0111; // x=112, y=22
        pixel_data[22][113] = 4'b0111; // x=113, y=22
        pixel_data[22][114] = 4'b0000; // x=114, y=22
        pixel_data[22][115] = 4'b0000; // x=115, y=22
        pixel_data[22][116] = 4'b0000; // x=116, y=22
        pixel_data[22][117] = 4'b0111; // x=117, y=22
        pixel_data[22][118] = 4'b0111; // x=118, y=22
        pixel_data[22][119] = 4'b0111; // x=119, y=22
        pixel_data[22][120] = 4'b0111; // x=120, y=22
        pixel_data[22][121] = 4'b0000; // x=121, y=22
        pixel_data[22][122] = 4'b0111; // x=122, y=22
        pixel_data[22][123] = 4'b0111; // x=123, y=22
        pixel_data[22][124] = 4'b0111; // x=124, y=22
        pixel_data[22][125] = 4'b0111; // x=125, y=22
        pixel_data[22][126] = 4'b0111; // x=126, y=22
        pixel_data[22][127] = 4'b0111; // x=127, y=22
        pixel_data[22][128] = 4'b0111; // x=128, y=22
        pixel_data[22][129] = 4'b0111; // x=129, y=22
        pixel_data[22][130] = 4'b0111; // x=130, y=22
        pixel_data[22][131] = 4'b0111; // x=131, y=22
        pixel_data[22][132] = 4'b0111; // x=132, y=22
        pixel_data[22][133] = 4'b0111; // x=133, y=22
        pixel_data[22][134] = 4'b0111; // x=134, y=22
        pixel_data[22][135] = 4'b0111; // x=135, y=22
        pixel_data[22][136] = 4'b0111; // x=136, y=22
        pixel_data[22][137] = 4'b0111; // x=137, y=22
        pixel_data[22][138] = 4'b0111; // x=138, y=22
        pixel_data[22][139] = 4'b0111; // x=139, y=22
        pixel_data[22][140] = 4'b0111; // x=140, y=22
        pixel_data[22][141] = 4'b0111; // x=141, y=22
        pixel_data[22][142] = 4'b0000; // x=142, y=22
        pixel_data[22][143] = 4'b0111; // x=143, y=22
        pixel_data[22][144] = 4'b0111; // x=144, y=22
        pixel_data[22][145] = 4'b0000; // x=145, y=22
        pixel_data[22][146] = 4'b0111; // x=146, y=22
        pixel_data[22][147] = 4'b0111; // x=147, y=22
        pixel_data[22][148] = 4'b0111; // x=148, y=22
        pixel_data[22][149] = 4'b0111; // x=149, y=22
        pixel_data[22][150] = 4'b0111; // x=150, y=22
        pixel_data[22][151] = 4'b0111; // x=151, y=22
        pixel_data[22][152] = 4'b0111; // x=152, y=22
        pixel_data[22][153] = 4'b0111; // x=153, y=22
        pixel_data[22][154] = 4'b0111; // x=154, y=22
        pixel_data[22][155] = 4'b0111; // x=155, y=22
        pixel_data[22][156] = 4'b0111; // x=156, y=22
        pixel_data[22][157] = 4'b0111; // x=157, y=22
        pixel_data[22][158] = 4'b0111; // x=158, y=22
        pixel_data[22][159] = 4'b0111; // x=159, y=22
        pixel_data[22][160] = 4'b0111; // x=160, y=22
        pixel_data[22][161] = 4'b0111; // x=161, y=22
        pixel_data[22][162] = 4'b0111; // x=162, y=22
        pixel_data[22][163] = 4'b0111; // x=163, y=22
        pixel_data[22][164] = 4'b0111; // x=164, y=22
        pixel_data[22][165] = 4'b0111; // x=165, y=22
        pixel_data[22][166] = 4'b0111; // x=166, y=22
        pixel_data[22][167] = 4'b0111; // x=167, y=22
        pixel_data[22][168] = 4'b0111; // x=168, y=22
        pixel_data[22][169] = 4'b0111; // x=169, y=22
        pixel_data[22][170] = 4'b0111; // x=170, y=22
        pixel_data[22][171] = 4'b0111; // x=171, y=22
        pixel_data[22][172] = 4'b0111; // x=172, y=22
        pixel_data[22][173] = 4'b0111; // x=173, y=22
        pixel_data[22][174] = 4'b0111; // x=174, y=22
        pixel_data[22][175] = 4'b0111; // x=175, y=22
        pixel_data[22][176] = 4'b0111; // x=176, y=22
        pixel_data[22][177] = 4'b0111; // x=177, y=22
        pixel_data[22][178] = 4'b0111; // x=178, y=22
        pixel_data[22][179] = 4'b0111; // x=179, y=22
        pixel_data[23][0] = 4'b0111; // x=0, y=23
        pixel_data[23][1] = 4'b0111; // x=1, y=23
        pixel_data[23][2] = 4'b0111; // x=2, y=23
        pixel_data[23][3] = 4'b0111; // x=3, y=23
        pixel_data[23][4] = 4'b0111; // x=4, y=23
        pixel_data[23][5] = 4'b0111; // x=5, y=23
        pixel_data[23][6] = 4'b0111; // x=6, y=23
        pixel_data[23][7] = 4'b0111; // x=7, y=23
        pixel_data[23][8] = 4'b0111; // x=8, y=23
        pixel_data[23][9] = 4'b0000; // x=9, y=23
        pixel_data[23][10] = 4'b1011; // x=10, y=23
        pixel_data[23][11] = 4'b1101; // x=11, y=23
        pixel_data[23][12] = 4'b1101; // x=12, y=23
        pixel_data[23][13] = 4'b0001; // x=13, y=23
        pixel_data[23][14] = 4'b1101; // x=14, y=23
        pixel_data[23][15] = 4'b1100; // x=15, y=23
        pixel_data[23][16] = 4'b0111; // x=16, y=23
        pixel_data[23][17] = 4'b0000; // x=17, y=23
        pixel_data[23][18] = 4'b0000; // x=18, y=23
        pixel_data[23][19] = 4'b0000; // x=19, y=23
        pixel_data[23][20] = 4'b0000; // x=20, y=23
        pixel_data[23][21] = 4'b0000; // x=21, y=23
        pixel_data[23][22] = 4'b0000; // x=22, y=23
        pixel_data[23][23] = 4'b0000; // x=23, y=23
        pixel_data[23][24] = 4'b0111; // x=24, y=23
        pixel_data[23][25] = 4'b0111; // x=25, y=23
        pixel_data[23][26] = 4'b1110; // x=26, y=23
        pixel_data[23][27] = 4'b1100; // x=27, y=23
        pixel_data[23][28] = 4'b1100; // x=28, y=23
        pixel_data[23][29] = 4'b1110; // x=29, y=23
        pixel_data[23][30] = 4'b0111; // x=30, y=23
        pixel_data[23][31] = 4'b0000; // x=31, y=23
        pixel_data[23][32] = 4'b0111; // x=32, y=23
        pixel_data[23][33] = 4'b0111; // x=33, y=23
        pixel_data[23][34] = 4'b0111; // x=34, y=23
        pixel_data[23][35] = 4'b0111; // x=35, y=23
        pixel_data[23][36] = 4'b0111; // x=36, y=23
        pixel_data[23][37] = 4'b0111; // x=37, y=23
        pixel_data[23][38] = 4'b0111; // x=38, y=23
        pixel_data[23][39] = 4'b0000; // x=39, y=23
        pixel_data[23][40] = 4'b0111; // x=40, y=23
        pixel_data[23][41] = 4'b0111; // x=41, y=23
        pixel_data[23][42] = 4'b0110; // x=42, y=23
        pixel_data[23][43] = 4'b1010; // x=43, y=23
        pixel_data[23][44] = 4'b1111; // x=44, y=23
        pixel_data[23][45] = 4'b1000; // x=45, y=23
        pixel_data[23][46] = 4'b0011; // x=46, y=23
        pixel_data[23][47] = 4'b0011; // x=47, y=23
        pixel_data[23][48] = 4'b1100; // x=48, y=23
        pixel_data[23][49] = 4'b1000; // x=49, y=23
        pixel_data[23][50] = 4'b0101; // x=50, y=23
        pixel_data[23][51] = 4'b1001; // x=51, y=23
        pixel_data[23][52] = 4'b1110; // x=52, y=23
        pixel_data[23][53] = 4'b0111; // x=53, y=23
        pixel_data[23][54] = 4'b0111; // x=54, y=23
        pixel_data[23][55] = 4'b0000; // x=55, y=23
        pixel_data[23][56] = 4'b0111; // x=56, y=23
        pixel_data[23][57] = 4'b0111; // x=57, y=23
        pixel_data[23][58] = 4'b0111; // x=58, y=23
        pixel_data[23][59] = 4'b0111; // x=59, y=23
        pixel_data[23][60] = 4'b0111; // x=60, y=23
        pixel_data[23][61] = 4'b0111; // x=61, y=23
        pixel_data[23][62] = 4'b0000; // x=62, y=23
        pixel_data[23][63] = 4'b0000; // x=63, y=23
        pixel_data[23][64] = 4'b0111; // x=64, y=23
        pixel_data[23][65] = 4'b0000; // x=65, y=23
        pixel_data[23][66] = 4'b0100; // x=66, y=23
        pixel_data[23][67] = 4'b0010; // x=67, y=23
        pixel_data[23][68] = 4'b1111; // x=68, y=23
        pixel_data[23][69] = 4'b1100; // x=69, y=23
        pixel_data[23][70] = 4'b0011; // x=70, y=23
        pixel_data[23][71] = 4'b0011; // x=71, y=23
        pixel_data[23][72] = 4'b1100; // x=72, y=23
        pixel_data[23][73] = 4'b1000; // x=73, y=23
        pixel_data[23][74] = 4'b0101; // x=74, y=23
        pixel_data[23][75] = 4'b0100; // x=75, y=23
        pixel_data[23][76] = 4'b1110; // x=76, y=23
        pixel_data[23][77] = 4'b0111; // x=77, y=23
        pixel_data[23][78] = 4'b0111; // x=78, y=23
        pixel_data[23][79] = 4'b0000; // x=79, y=23
        pixel_data[23][80] = 4'b0111; // x=80, y=23
        pixel_data[23][81] = 4'b0111; // x=81, y=23
        pixel_data[23][82] = 4'b0111; // x=82, y=23
        pixel_data[23][83] = 4'b0111; // x=83, y=23
        pixel_data[23][84] = 4'b0111; // x=84, y=23
        pixel_data[23][85] = 4'b0111; // x=85, y=23
        pixel_data[23][86] = 4'b0111; // x=86, y=23
        pixel_data[23][87] = 4'b1110; // x=87, y=23
        pixel_data[23][88] = 4'b0010; // x=88, y=23
        pixel_data[23][89] = 4'b0101; // x=89, y=23
        pixel_data[23][90] = 4'b0101; // x=90, y=23
        pixel_data[23][91] = 4'b0101; // x=91, y=23
        pixel_data[23][92] = 4'b0010; // x=92, y=23
        pixel_data[23][93] = 4'b0110; // x=93, y=23
        pixel_data[23][94] = 4'b0111; // x=94, y=23
        pixel_data[23][95] = 4'b0111; // x=95, y=23
        pixel_data[23][96] = 4'b1110; // x=96, y=23
        pixel_data[23][97] = 4'b0010; // x=97, y=23
        pixel_data[23][98] = 4'b1000; // x=98, y=23
        pixel_data[23][99] = 4'b0011; // x=99, y=23
        pixel_data[23][100] = 4'b0011; // x=100, y=23
        pixel_data[23][101] = 4'b1100; // x=101, y=23
        pixel_data[23][102] = 4'b1010; // x=102, y=23
        pixel_data[23][103] = 4'b0111; // x=103, y=23
        pixel_data[23][104] = 4'b0111; // x=104, y=23
        pixel_data[23][105] = 4'b0111; // x=105, y=23
        pixel_data[23][106] = 4'b0111; // x=106, y=23
        pixel_data[23][107] = 4'b0000; // x=107, y=23
        pixel_data[23][108] = 4'b0111; // x=108, y=23
        pixel_data[23][109] = 4'b0111; // x=109, y=23
        pixel_data[23][110] = 4'b0110; // x=110, y=23
        pixel_data[23][111] = 4'b1010; // x=111, y=23
        pixel_data[23][112] = 4'b1111; // x=112, y=23
        pixel_data[23][113] = 4'b1100; // x=113, y=23
        pixel_data[23][114] = 4'b0011; // x=114, y=23
        pixel_data[23][115] = 4'b0011; // x=115, y=23
        pixel_data[23][116] = 4'b0011; // x=116, y=23
        pixel_data[23][117] = 4'b1100; // x=117, y=23
        pixel_data[23][118] = 4'b0101; // x=118, y=23
        pixel_data[23][119] = 4'b1001; // x=119, y=23
        pixel_data[23][120] = 4'b0000; // x=120, y=23
        pixel_data[23][121] = 4'b0111; // x=121, y=23
        pixel_data[23][122] = 4'b0111; // x=122, y=23
        pixel_data[23][123] = 4'b0111; // x=123, y=23
        pixel_data[23][124] = 4'b0111; // x=124, y=23
        pixel_data[23][125] = 4'b0111; // x=125, y=23
        pixel_data[23][126] = 4'b0111; // x=126, y=23
        pixel_data[23][127] = 4'b0111; // x=127, y=23
        pixel_data[23][128] = 4'b0111; // x=128, y=23
        pixel_data[23][129] = 4'b0111; // x=129, y=23
        pixel_data[23][130] = 4'b0111; // x=130, y=23
        pixel_data[23][131] = 4'b0111; // x=131, y=23
        pixel_data[23][132] = 4'b0111; // x=132, y=23
        pixel_data[23][133] = 4'b0111; // x=133, y=23
        pixel_data[23][134] = 4'b0111; // x=134, y=23
        pixel_data[23][135] = 4'b0111; // x=135, y=23
        pixel_data[23][136] = 4'b0111; // x=136, y=23
        pixel_data[23][137] = 4'b0111; // x=137, y=23
        pixel_data[23][138] = 4'b0111; // x=138, y=23
        pixel_data[23][139] = 4'b0111; // x=139, y=23
        pixel_data[23][140] = 4'b0111; // x=140, y=23
        pixel_data[23][141] = 4'b0000; // x=141, y=23
        pixel_data[23][142] = 4'b0111; // x=142, y=23
        pixel_data[23][143] = 4'b0100; // x=143, y=23
        pixel_data[23][144] = 4'b1111; // x=144, y=23
        pixel_data[23][145] = 4'b1100; // x=145, y=23
        pixel_data[23][146] = 4'b1100; // x=146, y=23
        pixel_data[23][147] = 4'b0010; // x=147, y=23
        pixel_data[23][148] = 4'b0000; // x=148, y=23
        pixel_data[23][149] = 4'b0111; // x=149, y=23
        pixel_data[23][150] = 4'b0111; // x=150, y=23
        pixel_data[23][151] = 4'b0111; // x=151, y=23
        pixel_data[23][152] = 4'b0111; // x=152, y=23
        pixel_data[23][153] = 4'b0111; // x=153, y=23
        pixel_data[23][154] = 4'b0111; // x=154, y=23
        pixel_data[23][155] = 4'b0111; // x=155, y=23
        pixel_data[23][156] = 4'b0111; // x=156, y=23
        pixel_data[23][157] = 4'b0111; // x=157, y=23
        pixel_data[23][158] = 4'b0111; // x=158, y=23
        pixel_data[23][159] = 4'b0111; // x=159, y=23
        pixel_data[23][160] = 4'b0111; // x=160, y=23
        pixel_data[23][161] = 4'b0111; // x=161, y=23
        pixel_data[23][162] = 4'b0111; // x=162, y=23
        pixel_data[23][163] = 4'b0111; // x=163, y=23
        pixel_data[23][164] = 4'b0111; // x=164, y=23
        pixel_data[23][165] = 4'b0111; // x=165, y=23
        pixel_data[23][166] = 4'b0111; // x=166, y=23
        pixel_data[23][167] = 4'b0111; // x=167, y=23
        pixel_data[23][168] = 4'b0111; // x=168, y=23
        pixel_data[23][169] = 4'b0111; // x=169, y=23
        pixel_data[23][170] = 4'b0111; // x=170, y=23
        pixel_data[23][171] = 4'b0111; // x=171, y=23
        pixel_data[23][172] = 4'b0111; // x=172, y=23
        pixel_data[23][173] = 4'b0111; // x=173, y=23
        pixel_data[23][174] = 4'b0111; // x=174, y=23
        pixel_data[23][175] = 4'b0111; // x=175, y=23
        pixel_data[23][176] = 4'b0111; // x=176, y=23
        pixel_data[23][177] = 4'b0111; // x=177, y=23
        pixel_data[23][178] = 4'b0111; // x=178, y=23
        pixel_data[23][179] = 4'b0111; // x=179, y=23
        pixel_data[24][0] = 4'b0111; // x=0, y=24
        pixel_data[24][1] = 4'b0111; // x=1, y=24
        pixel_data[24][2] = 4'b0111; // x=2, y=24
        pixel_data[24][3] = 4'b0111; // x=3, y=24
        pixel_data[24][4] = 4'b0111; // x=4, y=24
        pixel_data[24][5] = 4'b0111; // x=5, y=24
        pixel_data[24][6] = 4'b0111; // x=6, y=24
        pixel_data[24][7] = 4'b0111; // x=7, y=24
        pixel_data[24][8] = 4'b0111; // x=8, y=24
        pixel_data[24][9] = 4'b0000; // x=9, y=24
        pixel_data[24][10] = 4'b1011; // x=10, y=24
        pixel_data[24][11] = 4'b1101; // x=11, y=24
        pixel_data[24][12] = 4'b0001; // x=12, y=24
        pixel_data[24][13] = 4'b0001; // x=13, y=24
        pixel_data[24][14] = 4'b1101; // x=14, y=24
        pixel_data[24][15] = 4'b0011; // x=15, y=24
        pixel_data[24][16] = 4'b0111; // x=16, y=24
        pixel_data[24][17] = 4'b0000; // x=17, y=24
        pixel_data[24][18] = 4'b0000; // x=18, y=24
        pixel_data[24][19] = 4'b0000; // x=19, y=24
        pixel_data[24][20] = 4'b0111; // x=20, y=24
        pixel_data[24][21] = 4'b0000; // x=21, y=24
        pixel_data[24][22] = 4'b0000; // x=22, y=24
        pixel_data[24][23] = 4'b0000; // x=23, y=24
        pixel_data[24][24] = 4'b0000; // x=24, y=24
        pixel_data[24][25] = 4'b0000; // x=25, y=24
        pixel_data[24][26] = 4'b0111; // x=26, y=24
        pixel_data[24][27] = 4'b0000; // x=27, y=24
        pixel_data[24][28] = 4'b0000; // x=28, y=24
        pixel_data[24][29] = 4'b0111; // x=29, y=24
        pixel_data[24][30] = 4'b0000; // x=30, y=24
        pixel_data[24][31] = 4'b0111; // x=31, y=24
        pixel_data[24][32] = 4'b0111; // x=32, y=24
        pixel_data[24][33] = 4'b0111; // x=33, y=24
        pixel_data[24][34] = 4'b0111; // x=34, y=24
        pixel_data[24][35] = 4'b0111; // x=35, y=24
        pixel_data[24][36] = 4'b0111; // x=36, y=24
        pixel_data[24][37] = 4'b0111; // x=37, y=24
        pixel_data[24][38] = 4'b0111; // x=38, y=24
        pixel_data[24][39] = 4'b0111; // x=39, y=24
        pixel_data[24][40] = 4'b0110; // x=40, y=24
        pixel_data[24][41] = 4'b1000; // x=41, y=24
        pixel_data[24][42] = 4'b1011; // x=42, y=24
        pixel_data[24][43] = 4'b1101; // x=43, y=24
        pixel_data[24][44] = 4'b1101; // x=44, y=24
        pixel_data[24][45] = 4'b1101; // x=45, y=24
        pixel_data[24][46] = 4'b1101; // x=46, y=24
        pixel_data[24][47] = 4'b1101; // x=47, y=24
        pixel_data[24][48] = 4'b1101; // x=48, y=24
        pixel_data[24][49] = 4'b1101; // x=49, y=24
        pixel_data[24][50] = 4'b1101; // x=50, y=24
        pixel_data[24][51] = 4'b1101; // x=51, y=24
        pixel_data[24][52] = 4'b1011; // x=52, y=24
        pixel_data[24][53] = 4'b0101; // x=53, y=24
        pixel_data[24][54] = 4'b0110; // x=54, y=24
        pixel_data[24][55] = 4'b0111; // x=55, y=24
        pixel_data[24][56] = 4'b0111; // x=56, y=24
        pixel_data[24][57] = 4'b0000; // x=57, y=24
        pixel_data[24][58] = 4'b0111; // x=58, y=24
        pixel_data[24][59] = 4'b0111; // x=59, y=24
        pixel_data[24][60] = 4'b0111; // x=60, y=24
        pixel_data[24][61] = 4'b0000; // x=61, y=24
        pixel_data[24][62] = 4'b0111; // x=62, y=24
        pixel_data[24][63] = 4'b0000; // x=63, y=24
        pixel_data[24][64] = 4'b1010; // x=64, y=24
        pixel_data[24][65] = 4'b0011; // x=65, y=24
        pixel_data[24][66] = 4'b0001; // x=66, y=24
        pixel_data[24][67] = 4'b1101; // x=67, y=24
        pixel_data[24][68] = 4'b1101; // x=68, y=24
        pixel_data[24][69] = 4'b1101; // x=69, y=24
        pixel_data[24][70] = 4'b1101; // x=70, y=24
        pixel_data[24][71] = 4'b1101; // x=71, y=24
        pixel_data[24][72] = 4'b1101; // x=72, y=24
        pixel_data[24][73] = 4'b1101; // x=73, y=24
        pixel_data[24][74] = 4'b1101; // x=74, y=24
        pixel_data[24][75] = 4'b1101; // x=75, y=24
        pixel_data[24][76] = 4'b0011; // x=76, y=24
        pixel_data[24][77] = 4'b0101; // x=77, y=24
        pixel_data[24][78] = 4'b1110; // x=78, y=24
        pixel_data[24][79] = 4'b0111; // x=79, y=24
        pixel_data[24][80] = 4'b0000; // x=80, y=24
        pixel_data[24][81] = 4'b0111; // x=81, y=24
        pixel_data[24][82] = 4'b0111; // x=82, y=24
        pixel_data[24][83] = 4'b0111; // x=83, y=24
        pixel_data[24][84] = 4'b0111; // x=84, y=24
        pixel_data[24][85] = 4'b0000; // x=85, y=24
        pixel_data[24][86] = 4'b0111; // x=86, y=24
        pixel_data[24][87] = 4'b0110; // x=87, y=24
        pixel_data[24][88] = 4'b1101; // x=88, y=24
        pixel_data[24][89] = 4'b1101; // x=89, y=24
        pixel_data[24][90] = 4'b1101; // x=90, y=24
        pixel_data[24][91] = 4'b1101; // x=91, y=24
        pixel_data[24][92] = 4'b1101; // x=92, y=24
        pixel_data[24][93] = 4'b0100; // x=93, y=24
        pixel_data[24][94] = 4'b0000; // x=94, y=24
        pixel_data[24][95] = 4'b0101; // x=95, y=24
        pixel_data[24][96] = 4'b1011; // x=96, y=24
        pixel_data[24][97] = 4'b1101; // x=97, y=24
        pixel_data[24][98] = 4'b1101; // x=98, y=24
        pixel_data[24][99] = 4'b1101; // x=99, y=24
        pixel_data[24][100] = 4'b1101; // x=100, y=24
        pixel_data[24][101] = 4'b1101; // x=101, y=24
        pixel_data[24][102] = 4'b1010; // x=102, y=24
        pixel_data[24][103] = 4'b0111; // x=103, y=24
        pixel_data[24][104] = 4'b0000; // x=104, y=24
        pixel_data[24][105] = 4'b0000; // x=105, y=24
        pixel_data[24][106] = 4'b0111; // x=106, y=24
        pixel_data[24][107] = 4'b0111; // x=107, y=24
        pixel_data[24][108] = 4'b0100; // x=108, y=24
        pixel_data[24][109] = 4'b1000; // x=109, y=24
        pixel_data[24][110] = 4'b0001; // x=110, y=24
        pixel_data[24][111] = 4'b1101; // x=111, y=24
        pixel_data[24][112] = 4'b1101; // x=112, y=24
        pixel_data[24][113] = 4'b1101; // x=113, y=24
        pixel_data[24][114] = 4'b1101; // x=114, y=24
        pixel_data[24][115] = 4'b1101; // x=115, y=24
        pixel_data[24][116] = 4'b1101; // x=116, y=24
        pixel_data[24][117] = 4'b1101; // x=117, y=24
        pixel_data[24][118] = 4'b1101; // x=118, y=24
        pixel_data[24][119] = 4'b1101; // x=119, y=24
        pixel_data[24][120] = 4'b0011; // x=120, y=24
        pixel_data[24][121] = 4'b1010; // x=121, y=24
        pixel_data[24][122] = 4'b0000; // x=122, y=24
        pixel_data[24][123] = 4'b0111; // x=123, y=24
        pixel_data[24][124] = 4'b0000; // x=124, y=24
        pixel_data[24][125] = 4'b0111; // x=125, y=24
        pixel_data[24][126] = 4'b0111; // x=126, y=24
        pixel_data[24][127] = 4'b0111; // x=127, y=24
        pixel_data[24][128] = 4'b0111; // x=128, y=24
        pixel_data[24][129] = 4'b0111; // x=129, y=24
        pixel_data[24][130] = 4'b0111; // x=130, y=24
        pixel_data[24][131] = 4'b0111; // x=131, y=24
        pixel_data[24][132] = 4'b0111; // x=132, y=24
        pixel_data[24][133] = 4'b0111; // x=133, y=24
        pixel_data[24][134] = 4'b0111; // x=134, y=24
        pixel_data[24][135] = 4'b0111; // x=135, y=24
        pixel_data[24][136] = 4'b0111; // x=136, y=24
        pixel_data[24][137] = 4'b0111; // x=137, y=24
        pixel_data[24][138] = 4'b0111; // x=138, y=24
        pixel_data[24][139] = 4'b0111; // x=139, y=24
        pixel_data[24][140] = 4'b0000; // x=140, y=24
        pixel_data[24][141] = 4'b0111; // x=141, y=24
        pixel_data[24][142] = 4'b0100; // x=142, y=24
        pixel_data[24][143] = 4'b0001; // x=143, y=24
        pixel_data[24][144] = 4'b1101; // x=144, y=24
        pixel_data[24][145] = 4'b1101; // x=145, y=24
        pixel_data[24][146] = 4'b1101; // x=146, y=24
        pixel_data[24][147] = 4'b1101; // x=147, y=24
        pixel_data[24][148] = 4'b0101; // x=148, y=24
        pixel_data[24][149] = 4'b0111; // x=149, y=24
        pixel_data[24][150] = 4'b0000; // x=150, y=24
        pixel_data[24][151] = 4'b0000; // x=151, y=24
        pixel_data[24][152] = 4'b0111; // x=152, y=24
        pixel_data[24][153] = 4'b0111; // x=153, y=24
        pixel_data[24][154] = 4'b0111; // x=154, y=24
        pixel_data[24][155] = 4'b0111; // x=155, y=24
        pixel_data[24][156] = 4'b0111; // x=156, y=24
        pixel_data[24][157] = 4'b0111; // x=157, y=24
        pixel_data[24][158] = 4'b0111; // x=158, y=24
        pixel_data[24][159] = 4'b0111; // x=159, y=24
        pixel_data[24][160] = 4'b0111; // x=160, y=24
        pixel_data[24][161] = 4'b0111; // x=161, y=24
        pixel_data[24][162] = 4'b0111; // x=162, y=24
        pixel_data[24][163] = 4'b0111; // x=163, y=24
        pixel_data[24][164] = 4'b0111; // x=164, y=24
        pixel_data[24][165] = 4'b0111; // x=165, y=24
        pixel_data[24][166] = 4'b0111; // x=166, y=24
        pixel_data[24][167] = 4'b0111; // x=167, y=24
        pixel_data[24][168] = 4'b0111; // x=168, y=24
        pixel_data[24][169] = 4'b0111; // x=169, y=24
        pixel_data[24][170] = 4'b0111; // x=170, y=24
        pixel_data[24][171] = 4'b0111; // x=171, y=24
        pixel_data[24][172] = 4'b0111; // x=172, y=24
        pixel_data[24][173] = 4'b0111; // x=173, y=24
        pixel_data[24][174] = 4'b0111; // x=174, y=24
        pixel_data[24][175] = 4'b0111; // x=175, y=24
        pixel_data[24][176] = 4'b0111; // x=176, y=24
        pixel_data[24][177] = 4'b0111; // x=177, y=24
        pixel_data[24][178] = 4'b0111; // x=178, y=24
        pixel_data[24][179] = 4'b0111; // x=179, y=24
        pixel_data[25][0] = 4'b0111; // x=0, y=25
        pixel_data[25][1] = 4'b0111; // x=1, y=25
        pixel_data[25][2] = 4'b0111; // x=2, y=25
        pixel_data[25][3] = 4'b0111; // x=3, y=25
        pixel_data[25][4] = 4'b0111; // x=4, y=25
        pixel_data[25][5] = 4'b0111; // x=5, y=25
        pixel_data[25][6] = 4'b0111; // x=6, y=25
        pixel_data[25][7] = 4'b0111; // x=7, y=25
        pixel_data[25][8] = 4'b0111; // x=8, y=25
        pixel_data[25][9] = 4'b0111; // x=9, y=25
        pixel_data[25][10] = 4'b0011; // x=10, y=25
        pixel_data[25][11] = 4'b1101; // x=11, y=25
        pixel_data[25][12] = 4'b0001; // x=12, y=25
        pixel_data[25][13] = 4'b1101; // x=13, y=25
        pixel_data[25][14] = 4'b1101; // x=14, y=25
        pixel_data[25][15] = 4'b1101; // x=15, y=25
        pixel_data[25][16] = 4'b0101; // x=16, y=25
        pixel_data[25][17] = 4'b0000; // x=17, y=25
        pixel_data[25][18] = 4'b0111; // x=18, y=25
        pixel_data[25][19] = 4'b0111; // x=19, y=25
        pixel_data[25][20] = 4'b0111; // x=20, y=25
        pixel_data[25][21] = 4'b0000; // x=21, y=25
        pixel_data[25][22] = 4'b0000; // x=22, y=25
        pixel_data[25][23] = 4'b0000; // x=23, y=25
        pixel_data[25][24] = 4'b0000; // x=24, y=25
        pixel_data[25][25] = 4'b0111; // x=25, y=25
        pixel_data[25][26] = 4'b0000; // x=26, y=25
        pixel_data[25][27] = 4'b0111; // x=27, y=25
        pixel_data[25][28] = 4'b0111; // x=28, y=25
        pixel_data[25][29] = 4'b0111; // x=29, y=25
        pixel_data[25][30] = 4'b0111; // x=30, y=25
        pixel_data[25][31] = 4'b0111; // x=31, y=25
        pixel_data[25][32] = 4'b0111; // x=32, y=25
        pixel_data[25][33] = 4'b0111; // x=33, y=25
        pixel_data[25][34] = 4'b0111; // x=34, y=25
        pixel_data[25][35] = 4'b0111; // x=35, y=25
        pixel_data[25][36] = 4'b0000; // x=36, y=25
        pixel_data[25][37] = 4'b0000; // x=37, y=25
        pixel_data[25][38] = 4'b0111; // x=38, y=25
        pixel_data[25][39] = 4'b0010; // x=39, y=25
        pixel_data[25][40] = 4'b0001; // x=40, y=25
        pixel_data[25][41] = 4'b1101; // x=41, y=25
        pixel_data[25][42] = 4'b1101; // x=42, y=25
        pixel_data[25][43] = 4'b0001; // x=43, y=25
        pixel_data[25][44] = 4'b1011; // x=44, y=25
        pixel_data[25][45] = 4'b0001; // x=45, y=25
        pixel_data[25][46] = 4'b1101; // x=46, y=25
        pixel_data[25][47] = 4'b1101; // x=47, y=25
        pixel_data[25][48] = 4'b1101; // x=48, y=25
        pixel_data[25][49] = 4'b0001; // x=49, y=25
        pixel_data[25][50] = 4'b0001; // x=50, y=25
        pixel_data[25][51] = 4'b0001; // x=51, y=25
        pixel_data[25][52] = 4'b1101; // x=52, y=25
        pixel_data[25][53] = 4'b1101; // x=53, y=25
        pixel_data[25][54] = 4'b0001; // x=54, y=25
        pixel_data[25][55] = 4'b1010; // x=55, y=25
        pixel_data[25][56] = 4'b0111; // x=56, y=25
        pixel_data[25][57] = 4'b0000; // x=57, y=25
        pixel_data[25][58] = 4'b0000; // x=58, y=25
        pixel_data[25][59] = 4'b0000; // x=59, y=25
        pixel_data[25][60] = 4'b0000; // x=60, y=25
        pixel_data[25][61] = 4'b0111; // x=61, y=25
        pixel_data[25][62] = 4'b0100; // x=62, y=25
        pixel_data[25][63] = 4'b1100; // x=63, y=25
        pixel_data[25][64] = 4'b1101; // x=64, y=25
        pixel_data[25][65] = 4'b1101; // x=65, y=25
        pixel_data[25][66] = 4'b0001; // x=66, y=25
        pixel_data[25][67] = 4'b0001; // x=67, y=25
        pixel_data[25][68] = 4'b0001; // x=68, y=25
        pixel_data[25][69] = 4'b1101; // x=69, y=25
        pixel_data[25][70] = 4'b1101; // x=70, y=25
        pixel_data[25][71] = 4'b1101; // x=71, y=25
        pixel_data[25][72] = 4'b1101; // x=72, y=25
        pixel_data[25][73] = 4'b0001; // x=73, y=25
        pixel_data[25][74] = 4'b0001; // x=74, y=25
        pixel_data[25][75] = 4'b0001; // x=75, y=25
        pixel_data[25][76] = 4'b1101; // x=76, y=25
        pixel_data[25][77] = 4'b1101; // x=77, y=25
        pixel_data[25][78] = 4'b0011; // x=78, y=25
        pixel_data[25][79] = 4'b1001; // x=79, y=25
        pixel_data[25][80] = 4'b0111; // x=80, y=25
        pixel_data[25][81] = 4'b0000; // x=81, y=25
        pixel_data[25][82] = 4'b0111; // x=82, y=25
        pixel_data[25][83] = 4'b0111; // x=83, y=25
        pixel_data[25][84] = 4'b0111; // x=84, y=25
        pixel_data[25][85] = 4'b0111; // x=85, y=25
        pixel_data[25][86] = 4'b0111; // x=86, y=25
        pixel_data[25][87] = 4'b0110; // x=87, y=25
        pixel_data[25][88] = 4'b1011; // x=88, y=25
        pixel_data[25][89] = 4'b0001; // x=89, y=25
        pixel_data[25][90] = 4'b0001; // x=90, y=25
        pixel_data[25][91] = 4'b0001; // x=91, y=25
        pixel_data[25][92] = 4'b0001; // x=92, y=25
        pixel_data[25][93] = 4'b1001; // x=93, y=25
        pixel_data[25][94] = 4'b1000; // x=94, y=25
        pixel_data[25][95] = 4'b1101; // x=95, y=25
        pixel_data[25][96] = 4'b1101; // x=96, y=25
        pixel_data[25][97] = 4'b0001; // x=97, y=25
        pixel_data[25][98] = 4'b0001; // x=98, y=25
        pixel_data[25][99] = 4'b0001; // x=99, y=25
        pixel_data[25][100] = 4'b0001; // x=100, y=25
        pixel_data[25][101] = 4'b1011; // x=101, y=25
        pixel_data[25][102] = 4'b0110; // x=102, y=25
        pixel_data[25][103] = 4'b0111; // x=103, y=25
        pixel_data[25][104] = 4'b0000; // x=104, y=25
        pixel_data[25][105] = 4'b0000; // x=105, y=25
        pixel_data[25][106] = 4'b0000; // x=106, y=25
        pixel_data[25][107] = 4'b0101; // x=107, y=25
        pixel_data[25][108] = 4'b1101; // x=108, y=25
        pixel_data[25][109] = 4'b1101; // x=109, y=25
        pixel_data[25][110] = 4'b1101; // x=110, y=25
        pixel_data[25][111] = 4'b0001; // x=111, y=25
        pixel_data[25][112] = 4'b0001; // x=112, y=25
        pixel_data[25][113] = 4'b1101; // x=113, y=25
        pixel_data[25][114] = 4'b1101; // x=114, y=25
        pixel_data[25][115] = 4'b1101; // x=115, y=25
        pixel_data[25][116] = 4'b1101; // x=116, y=25
        pixel_data[25][117] = 4'b0001; // x=117, y=25
        pixel_data[25][118] = 4'b0001; // x=118, y=25
        pixel_data[25][119] = 4'b0001; // x=119, y=25
        pixel_data[25][120] = 4'b1101; // x=120, y=25
        pixel_data[25][121] = 4'b1101; // x=121, y=25
        pixel_data[25][122] = 4'b1100; // x=122, y=25
        pixel_data[25][123] = 4'b1110; // x=123, y=25
        pixel_data[25][124] = 4'b0111; // x=124, y=25
        pixel_data[25][125] = 4'b0000; // x=125, y=25
        pixel_data[25][126] = 4'b0111; // x=126, y=25
        pixel_data[25][127] = 4'b0111; // x=127, y=25
        pixel_data[25][128] = 4'b0111; // x=128, y=25
        pixel_data[25][129] = 4'b0111; // x=129, y=25
        pixel_data[25][130] = 4'b0111; // x=130, y=25
        pixel_data[25][131] = 4'b0111; // x=131, y=25
        pixel_data[25][132] = 4'b0111; // x=132, y=25
        pixel_data[25][133] = 4'b0111; // x=133, y=25
        pixel_data[25][134] = 4'b0111; // x=134, y=25
        pixel_data[25][135] = 4'b0111; // x=135, y=25
        pixel_data[25][136] = 4'b0111; // x=136, y=25
        pixel_data[25][137] = 4'b0111; // x=137, y=25
        pixel_data[25][138] = 4'b0111; // x=138, y=25
        pixel_data[25][139] = 4'b0111; // x=139, y=25
        pixel_data[25][140] = 4'b0000; // x=140, y=25
        pixel_data[25][141] = 4'b0111; // x=141, y=25
        pixel_data[25][142] = 4'b0101; // x=142, y=25
        pixel_data[25][143] = 4'b1101; // x=143, y=25
        pixel_data[25][144] = 4'b0001; // x=144, y=25
        pixel_data[25][145] = 4'b1101; // x=145, y=25
        pixel_data[25][146] = 4'b0001; // x=146, y=25
        pixel_data[25][147] = 4'b1101; // x=147, y=25
        pixel_data[25][148] = 4'b0011; // x=148, y=25
        pixel_data[25][149] = 4'b0000; // x=149, y=25
        pixel_data[25][150] = 4'b0111; // x=150, y=25
        pixel_data[25][151] = 4'b0111; // x=151, y=25
        pixel_data[25][152] = 4'b0111; // x=152, y=25
        pixel_data[25][153] = 4'b0111; // x=153, y=25
        pixel_data[25][154] = 4'b0111; // x=154, y=25
        pixel_data[25][155] = 4'b0111; // x=155, y=25
        pixel_data[25][156] = 4'b0111; // x=156, y=25
        pixel_data[25][157] = 4'b0111; // x=157, y=25
        pixel_data[25][158] = 4'b0111; // x=158, y=25
        pixel_data[25][159] = 4'b0111; // x=159, y=25
        pixel_data[25][160] = 4'b0111; // x=160, y=25
        pixel_data[25][161] = 4'b0111; // x=161, y=25
        pixel_data[25][162] = 4'b0111; // x=162, y=25
        pixel_data[25][163] = 4'b0111; // x=163, y=25
        pixel_data[25][164] = 4'b0111; // x=164, y=25
        pixel_data[25][165] = 4'b0111; // x=165, y=25
        pixel_data[25][166] = 4'b0111; // x=166, y=25
        pixel_data[25][167] = 4'b0111; // x=167, y=25
        pixel_data[25][168] = 4'b0111; // x=168, y=25
        pixel_data[25][169] = 4'b0111; // x=169, y=25
        pixel_data[25][170] = 4'b0111; // x=170, y=25
        pixel_data[25][171] = 4'b0111; // x=171, y=25
        pixel_data[25][172] = 4'b0111; // x=172, y=25
        pixel_data[25][173] = 4'b0111; // x=173, y=25
        pixel_data[25][174] = 4'b0111; // x=174, y=25
        pixel_data[25][175] = 4'b0111; // x=175, y=25
        pixel_data[25][176] = 4'b0111; // x=176, y=25
        pixel_data[25][177] = 4'b0111; // x=177, y=25
        pixel_data[25][178] = 4'b0111; // x=178, y=25
        pixel_data[25][179] = 4'b0111; // x=179, y=25
        pixel_data[26][0] = 4'b0111; // x=0, y=26
        pixel_data[26][1] = 4'b0111; // x=1, y=26
        pixel_data[26][2] = 4'b0111; // x=2, y=26
        pixel_data[26][3] = 4'b0111; // x=3, y=26
        pixel_data[26][4] = 4'b0111; // x=4, y=26
        pixel_data[26][5] = 4'b0111; // x=5, y=26
        pixel_data[26][6] = 4'b0111; // x=6, y=26
        pixel_data[26][7] = 4'b0111; // x=7, y=26
        pixel_data[26][8] = 4'b0111; // x=8, y=26
        pixel_data[26][9] = 4'b0111; // x=9, y=26
        pixel_data[26][10] = 4'b0010; // x=10, y=26
        pixel_data[26][11] = 4'b1101; // x=11, y=26
        pixel_data[26][12] = 4'b0001; // x=12, y=26
        pixel_data[26][13] = 4'b1101; // x=13, y=26
        pixel_data[26][14] = 4'b0001; // x=14, y=26
        pixel_data[26][15] = 4'b0001; // x=15, y=26
        pixel_data[26][16] = 4'b1101; // x=16, y=26
        pixel_data[26][17] = 4'b0011; // x=17, y=26
        pixel_data[26][18] = 4'b0010; // x=18, y=26
        pixel_data[26][19] = 4'b0110; // x=19, y=26
        pixel_data[26][20] = 4'b1110; // x=20, y=26
        pixel_data[26][21] = 4'b0111; // x=21, y=26
        pixel_data[26][22] = 4'b0111; // x=22, y=26
        pixel_data[26][23] = 4'b0111; // x=23, y=26
        pixel_data[26][24] = 4'b0111; // x=24, y=26
        pixel_data[26][25] = 4'b0000; // x=25, y=26
        pixel_data[26][26] = 4'b0000; // x=26, y=26
        pixel_data[26][27] = 4'b0000; // x=27, y=26
        pixel_data[26][28] = 4'b0111; // x=28, y=26
        pixel_data[26][29] = 4'b0111; // x=29, y=26
        pixel_data[26][30] = 4'b0111; // x=30, y=26
        pixel_data[26][31] = 4'b0111; // x=31, y=26
        pixel_data[26][32] = 4'b0111; // x=32, y=26
        pixel_data[26][33] = 4'b0111; // x=33, y=26
        pixel_data[26][34] = 4'b0111; // x=34, y=26
        pixel_data[26][35] = 4'b0111; // x=35, y=26
        pixel_data[26][36] = 4'b0000; // x=36, y=26
        pixel_data[26][37] = 4'b0111; // x=37, y=26
        pixel_data[26][38] = 4'b0101; // x=38, y=26
        pixel_data[26][39] = 4'b1101; // x=39, y=26
        pixel_data[26][40] = 4'b0001; // x=40, y=26
        pixel_data[26][41] = 4'b0001; // x=41, y=26
        pixel_data[26][42] = 4'b0001; // x=42, y=26
        pixel_data[26][43] = 4'b1101; // x=43, y=26
        pixel_data[26][44] = 4'b1101; // x=44, y=26
        pixel_data[26][45] = 4'b0001; // x=45, y=26
        pixel_data[26][46] = 4'b1011; // x=46, y=26
        pixel_data[26][47] = 4'b0011; // x=47, y=26
        pixel_data[26][48] = 4'b1011; // x=48, y=26
        pixel_data[26][49] = 4'b0001; // x=49, y=26
        pixel_data[26][50] = 4'b1101; // x=50, y=26
        pixel_data[26][51] = 4'b1101; // x=51, y=26
        pixel_data[26][52] = 4'b0001; // x=52, y=26
        pixel_data[26][53] = 4'b0001; // x=53, y=26
        pixel_data[26][54] = 4'b0001; // x=54, y=26
        pixel_data[26][55] = 4'b1101; // x=55, y=26
        pixel_data[26][56] = 4'b1010; // x=56, y=26
        pixel_data[26][57] = 4'b0111; // x=57, y=26
        pixel_data[26][58] = 4'b0000; // x=58, y=26
        pixel_data[26][59] = 4'b0000; // x=59, y=26
        pixel_data[26][60] = 4'b0111; // x=60, y=26
        pixel_data[26][61] = 4'b0100; // x=61, y=26
        pixel_data[26][62] = 4'b1011; // x=62, y=26
        pixel_data[26][63] = 4'b1101; // x=63, y=26
        pixel_data[26][64] = 4'b0001; // x=64, y=26
        pixel_data[26][65] = 4'b0001; // x=65, y=26
        pixel_data[26][66] = 4'b0001; // x=66, y=26
        pixel_data[26][67] = 4'b1101; // x=67, y=26
        pixel_data[26][68] = 4'b1101; // x=68, y=26
        pixel_data[26][69] = 4'b1011; // x=69, y=26
        pixel_data[26][70] = 4'b0011; // x=70, y=26
        pixel_data[26][71] = 4'b0011; // x=71, y=26
        pixel_data[26][72] = 4'b1011; // x=72, y=26
        pixel_data[26][73] = 4'b1101; // x=73, y=26
        pixel_data[26][74] = 4'b1101; // x=74, y=26
        pixel_data[26][75] = 4'b1101; // x=75, y=26
        pixel_data[26][76] = 4'b0001; // x=76, y=26
        pixel_data[26][77] = 4'b0001; // x=77, y=26
        pixel_data[26][78] = 4'b1101; // x=78, y=26
        pixel_data[26][79] = 4'b1101; // x=79, y=26
        pixel_data[26][80] = 4'b1010; // x=80, y=26
        pixel_data[26][81] = 4'b0111; // x=81, y=26
        pixel_data[26][82] = 4'b0000; // x=82, y=26
        pixel_data[26][83] = 4'b0111; // x=83, y=26
        pixel_data[26][84] = 4'b0111; // x=84, y=26
        pixel_data[26][85] = 4'b0000; // x=85, y=26
        pixel_data[26][86] = 4'b0111; // x=86, y=26
        pixel_data[26][87] = 4'b0110; // x=87, y=26
        pixel_data[26][88] = 4'b1011; // x=88, y=26
        pixel_data[26][89] = 4'b1101; // x=89, y=26
        pixel_data[26][90] = 4'b1101; // x=90, y=26
        pixel_data[26][91] = 4'b1101; // x=91, y=26
        pixel_data[26][92] = 4'b0001; // x=92, y=26
        pixel_data[26][93] = 4'b1011; // x=93, y=26
        pixel_data[26][94] = 4'b1101; // x=94, y=26
        pixel_data[26][95] = 4'b0001; // x=95, y=26
        pixel_data[26][96] = 4'b1101; // x=96, y=26
        pixel_data[26][97] = 4'b1101; // x=97, y=26
        pixel_data[26][98] = 4'b1101; // x=98, y=26
        pixel_data[26][99] = 4'b1101; // x=99, y=26
        pixel_data[26][100] = 4'b1101; // x=100, y=26
        pixel_data[26][101] = 4'b1100; // x=101, y=26
        pixel_data[26][102] = 4'b0111; // x=102, y=26
        pixel_data[26][103] = 4'b0000; // x=103, y=26
        pixel_data[26][104] = 4'b0000; // x=104, y=26
        pixel_data[26][105] = 4'b0000; // x=105, y=26
        pixel_data[26][106] = 4'b1111; // x=106, y=26
        pixel_data[26][107] = 4'b1101; // x=107, y=26
        pixel_data[26][108] = 4'b1101; // x=108, y=26
        pixel_data[26][109] = 4'b0001; // x=109, y=26
        pixel_data[26][110] = 4'b0001; // x=110, y=26
        pixel_data[26][111] = 4'b1101; // x=111, y=26
        pixel_data[26][112] = 4'b1101; // x=112, y=26
        pixel_data[26][113] = 4'b1011; // x=113, y=26
        pixel_data[26][114] = 4'b0011; // x=114, y=26
        pixel_data[26][115] = 4'b1100; // x=115, y=26
        pixel_data[26][116] = 4'b0011; // x=116, y=26
        pixel_data[26][117] = 4'b0001; // x=117, y=26
        pixel_data[26][118] = 4'b1101; // x=118, y=26
        pixel_data[26][119] = 4'b1101; // x=119, y=26
        pixel_data[26][120] = 4'b0001; // x=120, y=26
        pixel_data[26][121] = 4'b0001; // x=121, y=26
        pixel_data[26][122] = 4'b1101; // x=122, y=26
        pixel_data[26][123] = 4'b0011; // x=123, y=26
        pixel_data[26][124] = 4'b1110; // x=124, y=26
        pixel_data[26][125] = 4'b0000; // x=125, y=26
        pixel_data[26][126] = 4'b0111; // x=126, y=26
        pixel_data[26][127] = 4'b0111; // x=127, y=26
        pixel_data[26][128] = 4'b0111; // x=128, y=26
        pixel_data[26][129] = 4'b0111; // x=129, y=26
        pixel_data[26][130] = 4'b0111; // x=130, y=26
        pixel_data[26][131] = 4'b0111; // x=131, y=26
        pixel_data[26][132] = 4'b0111; // x=132, y=26
        pixel_data[26][133] = 4'b0111; // x=133, y=26
        pixel_data[26][134] = 4'b0111; // x=134, y=26
        pixel_data[26][135] = 4'b0111; // x=135, y=26
        pixel_data[26][136] = 4'b0111; // x=136, y=26
        pixel_data[26][137] = 4'b0111; // x=137, y=26
        pixel_data[26][138] = 4'b0111; // x=138, y=26
        pixel_data[26][139] = 4'b0111; // x=139, y=26
        pixel_data[26][140] = 4'b0000; // x=140, y=26
        pixel_data[26][141] = 4'b0111; // x=141, y=26
        pixel_data[26][142] = 4'b0010; // x=142, y=26
        pixel_data[26][143] = 4'b1101; // x=143, y=26
        pixel_data[26][144] = 4'b0001; // x=144, y=26
        pixel_data[26][145] = 4'b1101; // x=145, y=26
        pixel_data[26][146] = 4'b0001; // x=146, y=26
        pixel_data[26][147] = 4'b1101; // x=147, y=26
        pixel_data[26][148] = 4'b1100; // x=148, y=26
        pixel_data[26][149] = 4'b0000; // x=149, y=26
        pixel_data[26][150] = 4'b0111; // x=150, y=26
        pixel_data[26][151] = 4'b0111; // x=151, y=26
        pixel_data[26][152] = 4'b0111; // x=152, y=26
        pixel_data[26][153] = 4'b0111; // x=153, y=26
        pixel_data[26][154] = 4'b0111; // x=154, y=26
        pixel_data[26][155] = 4'b0111; // x=155, y=26
        pixel_data[26][156] = 4'b0111; // x=156, y=26
        pixel_data[26][157] = 4'b0111; // x=157, y=26
        pixel_data[26][158] = 4'b0111; // x=158, y=26
        pixel_data[26][159] = 4'b0111; // x=159, y=26
        pixel_data[26][160] = 4'b0111; // x=160, y=26
        pixel_data[26][161] = 4'b0111; // x=161, y=26
        pixel_data[26][162] = 4'b0111; // x=162, y=26
        pixel_data[26][163] = 4'b0111; // x=163, y=26
        pixel_data[26][164] = 4'b0111; // x=164, y=26
        pixel_data[26][165] = 4'b0111; // x=165, y=26
        pixel_data[26][166] = 4'b0111; // x=166, y=26
        pixel_data[26][167] = 4'b0111; // x=167, y=26
        pixel_data[26][168] = 4'b0111; // x=168, y=26
        pixel_data[26][169] = 4'b0111; // x=169, y=26
        pixel_data[26][170] = 4'b0111; // x=170, y=26
        pixel_data[26][171] = 4'b0111; // x=171, y=26
        pixel_data[26][172] = 4'b0111; // x=172, y=26
        pixel_data[26][173] = 4'b0111; // x=173, y=26
        pixel_data[26][174] = 4'b0111; // x=174, y=26
        pixel_data[26][175] = 4'b0111; // x=175, y=26
        pixel_data[26][176] = 4'b0111; // x=176, y=26
        pixel_data[26][177] = 4'b0111; // x=177, y=26
        pixel_data[26][178] = 4'b0111; // x=178, y=26
        pixel_data[26][179] = 4'b0111; // x=179, y=26
        pixel_data[27][0] = 4'b0111; // x=0, y=27
        pixel_data[27][1] = 4'b0111; // x=1, y=27
        pixel_data[27][2] = 4'b0111; // x=2, y=27
        pixel_data[27][3] = 4'b0111; // x=3, y=27
        pixel_data[27][4] = 4'b0111; // x=4, y=27
        pixel_data[27][5] = 4'b0111; // x=5, y=27
        pixel_data[27][6] = 4'b0111; // x=6, y=27
        pixel_data[27][7] = 4'b0111; // x=7, y=27
        pixel_data[27][8] = 4'b0111; // x=8, y=27
        pixel_data[27][9] = 4'b0111; // x=9, y=27
        pixel_data[27][10] = 4'b1110; // x=10, y=27
        pixel_data[27][11] = 4'b0011; // x=11, y=27
        pixel_data[27][12] = 4'b1101; // x=12, y=27
        pixel_data[27][13] = 4'b0001; // x=13, y=27
        pixel_data[27][14] = 4'b0001; // x=14, y=27
        pixel_data[27][15] = 4'b0001; // x=15, y=27
        pixel_data[27][16] = 4'b0001; // x=16, y=27
        pixel_data[27][17] = 4'b1101; // x=17, y=27
        pixel_data[27][18] = 4'b1101; // x=18, y=27
        pixel_data[27][19] = 4'b1101; // x=19, y=27
        pixel_data[27][20] = 4'b0011; // x=20, y=27
        pixel_data[27][21] = 4'b1000; // x=21, y=27
        pixel_data[27][22] = 4'b0101; // x=22, y=27
        pixel_data[27][23] = 4'b1001; // x=23, y=27
        pixel_data[27][24] = 4'b0110; // x=24, y=27
        pixel_data[27][25] = 4'b0111; // x=25, y=27
        pixel_data[27][26] = 4'b0111; // x=26, y=27
        pixel_data[27][27] = 4'b0111; // x=27, y=27
        pixel_data[27][28] = 4'b0000; // x=28, y=27
        pixel_data[27][29] = 4'b0111; // x=29, y=27
        pixel_data[27][30] = 4'b0111; // x=30, y=27
        pixel_data[27][31] = 4'b0111; // x=31, y=27
        pixel_data[27][32] = 4'b0111; // x=32, y=27
        pixel_data[27][33] = 4'b0111; // x=33, y=27
        pixel_data[27][34] = 4'b0111; // x=34, y=27
        pixel_data[27][35] = 4'b0111; // x=35, y=27
        pixel_data[27][36] = 4'b0111; // x=36, y=27
        pixel_data[27][37] = 4'b0010; // x=37, y=27
        pixel_data[27][38] = 4'b1101; // x=38, y=27
        pixel_data[27][39] = 4'b0001; // x=39, y=27
        pixel_data[27][40] = 4'b0001; // x=40, y=27
        pixel_data[27][41] = 4'b0001; // x=41, y=27
        pixel_data[27][42] = 4'b1101; // x=42, y=27
        pixel_data[27][43] = 4'b1011; // x=43, y=27
        pixel_data[27][44] = 4'b0010; // x=44, y=27
        pixel_data[27][45] = 4'b0110; // x=45, y=27
        pixel_data[27][46] = 4'b0000; // x=46, y=27
        pixel_data[27][47] = 4'b0000; // x=47, y=27
        pixel_data[27][48] = 4'b0000; // x=48, y=27
        pixel_data[27][49] = 4'b0110; // x=49, y=27
        pixel_data[27][50] = 4'b1010; // x=50, y=27
        pixel_data[27][51] = 4'b0011; // x=51, y=27
        pixel_data[27][52] = 4'b1101; // x=52, y=27
        pixel_data[27][53] = 4'b1101; // x=53, y=27
        pixel_data[27][54] = 4'b1101; // x=54, y=27
        pixel_data[27][55] = 4'b1111; // x=55, y=27
        pixel_data[27][56] = 4'b1110; // x=56, y=27
        pixel_data[27][57] = 4'b0000; // x=57, y=27
        pixel_data[27][58] = 4'b0000; // x=58, y=27
        pixel_data[27][59] = 4'b0111; // x=59, y=27
        pixel_data[27][60] = 4'b0110; // x=60, y=27
        pixel_data[27][61] = 4'b1011; // x=61, y=27
        pixel_data[27][62] = 4'b1101; // x=62, y=27
        pixel_data[27][63] = 4'b0001; // x=63, y=27
        pixel_data[27][64] = 4'b0001; // x=64, y=27
        pixel_data[27][65] = 4'b1101; // x=65, y=27
        pixel_data[27][66] = 4'b1101; // x=66, y=27
        pixel_data[27][67] = 4'b1000; // x=67, y=27
        pixel_data[27][68] = 4'b1001; // x=68, y=27
        pixel_data[27][69] = 4'b1110; // x=69, y=27
        pixel_data[27][70] = 4'b0000; // x=70, y=27
        pixel_data[27][71] = 4'b0111; // x=71, y=27
        pixel_data[27][72] = 4'b1110; // x=72, y=27
        pixel_data[27][73] = 4'b0100; // x=73, y=27
        pixel_data[27][74] = 4'b1111; // x=74, y=27
        pixel_data[27][75] = 4'b1101; // x=75, y=27
        pixel_data[27][76] = 4'b1101; // x=76, y=27
        pixel_data[27][77] = 4'b0001; // x=77, y=27
        pixel_data[27][78] = 4'b0001; // x=78, y=27
        pixel_data[27][79] = 4'b0001; // x=79, y=27
        pixel_data[27][80] = 4'b1101; // x=80, y=27
        pixel_data[27][81] = 4'b1001; // x=81, y=27
        pixel_data[27][82] = 4'b0111; // x=82, y=27
        pixel_data[27][83] = 4'b0000; // x=83, y=27
        pixel_data[27][84] = 4'b0000; // x=84, y=27
        pixel_data[27][85] = 4'b0111; // x=85, y=27
        pixel_data[27][86] = 4'b0111; // x=86, y=27
        pixel_data[27][87] = 4'b0110; // x=87, y=27
        pixel_data[27][88] = 4'b1011; // x=88, y=27
        pixel_data[27][89] = 4'b1101; // x=89, y=27
        pixel_data[27][90] = 4'b1101; // x=90, y=27
        pixel_data[27][91] = 4'b1101; // x=91, y=27
        pixel_data[27][92] = 4'b1101; // x=92, y=27
        pixel_data[27][93] = 4'b1101; // x=93, y=27
        pixel_data[27][94] = 4'b1101; // x=94, y=27
        pixel_data[27][95] = 4'b1101; // x=95, y=27
        pixel_data[27][96] = 4'b1011; // x=96, y=27
        pixel_data[27][97] = 4'b1100; // x=97, y=27
        pixel_data[27][98] = 4'b1111; // x=98, y=27
        pixel_data[27][99] = 4'b1111; // x=99, y=27
        pixel_data[27][100] = 4'b0011; // x=100, y=27
        pixel_data[27][101] = 4'b1010; // x=101, y=27
        pixel_data[27][102] = 4'b0111; // x=102, y=27
        pixel_data[27][103] = 4'b0000; // x=103, y=27
        pixel_data[27][104] = 4'b0111; // x=104, y=27
        pixel_data[27][105] = 4'b0101; // x=105, y=27
        pixel_data[27][106] = 4'b1101; // x=106, y=27
        pixel_data[27][107] = 4'b0001; // x=107, y=27
        pixel_data[27][108] = 4'b0001; // x=108, y=27
        pixel_data[27][109] = 4'b0001; // x=109, y=27
        pixel_data[27][110] = 4'b0001; // x=110, y=27
        pixel_data[27][111] = 4'b1111; // x=111, y=27
        pixel_data[27][112] = 4'b0100; // x=112, y=27
        pixel_data[27][113] = 4'b1110; // x=113, y=27
        pixel_data[27][114] = 4'b0000; // x=114, y=27
        pixel_data[27][115] = 4'b0111; // x=115, y=27
        pixel_data[27][116] = 4'b0000; // x=116, y=27
        pixel_data[27][117] = 4'b0110; // x=117, y=27
        pixel_data[27][118] = 4'b0101; // x=118, y=27
        pixel_data[27][119] = 4'b0001; // x=119, y=27
        pixel_data[27][120] = 4'b0001; // x=120, y=27
        pixel_data[27][121] = 4'b0001; // x=121, y=27
        pixel_data[27][122] = 4'b0001; // x=122, y=27
        pixel_data[27][123] = 4'b1101; // x=123, y=27
        pixel_data[27][124] = 4'b1000; // x=124, y=27
        pixel_data[27][125] = 4'b0111; // x=125, y=27
        pixel_data[27][126] = 4'b0111; // x=126, y=27
        pixel_data[27][127] = 4'b0111; // x=127, y=27
        pixel_data[27][128] = 4'b0111; // x=128, y=27
        pixel_data[27][129] = 4'b0111; // x=129, y=27
        pixel_data[27][130] = 4'b0111; // x=130, y=27
        pixel_data[27][131] = 4'b0111; // x=131, y=27
        pixel_data[27][132] = 4'b0111; // x=132, y=27
        pixel_data[27][133] = 4'b0111; // x=133, y=27
        pixel_data[27][134] = 4'b0111; // x=134, y=27
        pixel_data[27][135] = 4'b0111; // x=135, y=27
        pixel_data[27][136] = 4'b0111; // x=136, y=27
        pixel_data[27][137] = 4'b0111; // x=137, y=27
        pixel_data[27][138] = 4'b0111; // x=138, y=27
        pixel_data[27][139] = 4'b0111; // x=139, y=27
        pixel_data[27][140] = 4'b0000; // x=140, y=27
        pixel_data[27][141] = 4'b0111; // x=141, y=27
        pixel_data[27][142] = 4'b0110; // x=142, y=27
        pixel_data[27][143] = 4'b0011; // x=143, y=27
        pixel_data[27][144] = 4'b1101; // x=144, y=27
        pixel_data[27][145] = 4'b1101; // x=145, y=27
        pixel_data[27][146] = 4'b1101; // x=146, y=27
        pixel_data[27][147] = 4'b1011; // x=147, y=27
        pixel_data[27][148] = 4'b1001; // x=148, y=27
        pixel_data[27][149] = 4'b0111; // x=149, y=27
        pixel_data[27][150] = 4'b0000; // x=150, y=27
        pixel_data[27][151] = 4'b0000; // x=151, y=27
        pixel_data[27][152] = 4'b0111; // x=152, y=27
        pixel_data[27][153] = 4'b0111; // x=153, y=27
        pixel_data[27][154] = 4'b0111; // x=154, y=27
        pixel_data[27][155] = 4'b0111; // x=155, y=27
        pixel_data[27][156] = 4'b0111; // x=156, y=27
        pixel_data[27][157] = 4'b0111; // x=157, y=27
        pixel_data[27][158] = 4'b0111; // x=158, y=27
        pixel_data[27][159] = 4'b0111; // x=159, y=27
        pixel_data[27][160] = 4'b0111; // x=160, y=27
        pixel_data[27][161] = 4'b0111; // x=161, y=27
        pixel_data[27][162] = 4'b0111; // x=162, y=27
        pixel_data[27][163] = 4'b0111; // x=163, y=27
        pixel_data[27][164] = 4'b0111; // x=164, y=27
        pixel_data[27][165] = 4'b0111; // x=165, y=27
        pixel_data[27][166] = 4'b0111; // x=166, y=27
        pixel_data[27][167] = 4'b0111; // x=167, y=27
        pixel_data[27][168] = 4'b0111; // x=168, y=27
        pixel_data[27][169] = 4'b0111; // x=169, y=27
        pixel_data[27][170] = 4'b0111; // x=170, y=27
        pixel_data[27][171] = 4'b0111; // x=171, y=27
        pixel_data[27][172] = 4'b0111; // x=172, y=27
        pixel_data[27][173] = 4'b0111; // x=173, y=27
        pixel_data[27][174] = 4'b0111; // x=174, y=27
        pixel_data[27][175] = 4'b0111; // x=175, y=27
        pixel_data[27][176] = 4'b0111; // x=176, y=27
        pixel_data[27][177] = 4'b0111; // x=177, y=27
        pixel_data[27][178] = 4'b0111; // x=178, y=27
        pixel_data[27][179] = 4'b0111; // x=179, y=27
        pixel_data[28][0] = 4'b0111; // x=0, y=28
        pixel_data[28][1] = 4'b0111; // x=1, y=28
        pixel_data[28][2] = 4'b0111; // x=2, y=28
        pixel_data[28][3] = 4'b0111; // x=3, y=28
        pixel_data[28][4] = 4'b0111; // x=4, y=28
        pixel_data[28][5] = 4'b0111; // x=5, y=28
        pixel_data[28][6] = 4'b0111; // x=6, y=28
        pixel_data[28][7] = 4'b0111; // x=7, y=28
        pixel_data[28][8] = 4'b0111; // x=8, y=28
        pixel_data[28][9] = 4'b0000; // x=9, y=28
        pixel_data[28][10] = 4'b0111; // x=10, y=28
        pixel_data[28][11] = 4'b0110; // x=11, y=28
        pixel_data[28][12] = 4'b0011; // x=12, y=28
        pixel_data[28][13] = 4'b1101; // x=13, y=28
        pixel_data[28][14] = 4'b1101; // x=14, y=28
        pixel_data[28][15] = 4'b0001; // x=15, y=28
        pixel_data[28][16] = 4'b0001; // x=16, y=28
        pixel_data[28][17] = 4'b0001; // x=17, y=28
        pixel_data[28][18] = 4'b0001; // x=18, y=28
        pixel_data[28][19] = 4'b1101; // x=19, y=28
        pixel_data[28][20] = 4'b1101; // x=20, y=28
        pixel_data[28][21] = 4'b1101; // x=21, y=28
        pixel_data[28][22] = 4'b1101; // x=22, y=28
        pixel_data[28][23] = 4'b1101; // x=23, y=28
        pixel_data[28][24] = 4'b0001; // x=24, y=28
        pixel_data[28][25] = 4'b1100; // x=25, y=28
        pixel_data[28][26] = 4'b0010; // x=26, y=28
        pixel_data[28][27] = 4'b0110; // x=27, y=28
        pixel_data[28][28] = 4'b0111; // x=28, y=28
        pixel_data[28][29] = 4'b0111; // x=29, y=28
        pixel_data[28][30] = 4'b0000; // x=30, y=28
        pixel_data[28][31] = 4'b0111; // x=31, y=28
        pixel_data[28][32] = 4'b0111; // x=32, y=28
        pixel_data[28][33] = 4'b0111; // x=33, y=28
        pixel_data[28][34] = 4'b0111; // x=34, y=28
        pixel_data[28][35] = 4'b0111; // x=35, y=28
        pixel_data[28][36] = 4'b0110; // x=36, y=28
        pixel_data[28][37] = 4'b0001; // x=37, y=28
        pixel_data[28][38] = 4'b0001; // x=38, y=28
        pixel_data[28][39] = 4'b0001; // x=39, y=28
        pixel_data[28][40] = 4'b0001; // x=40, y=28
        pixel_data[28][41] = 4'b1101; // x=41, y=28
        pixel_data[28][42] = 4'b1100; // x=42, y=28
        pixel_data[28][43] = 4'b0110; // x=43, y=28
        pixel_data[28][44] = 4'b0111; // x=44, y=28
        pixel_data[28][45] = 4'b0111; // x=45, y=28
        pixel_data[28][46] = 4'b0111; // x=46, y=28
        pixel_data[28][47] = 4'b0111; // x=47, y=28
        pixel_data[28][48] = 4'b0111; // x=48, y=28
        pixel_data[28][49] = 4'b0111; // x=49, y=28
        pixel_data[28][50] = 4'b0111; // x=50, y=28
        pixel_data[28][51] = 4'b0000; // x=51, y=28
        pixel_data[28][52] = 4'b0010; // x=52, y=28
        pixel_data[28][53] = 4'b0001; // x=53, y=28
        pixel_data[28][54] = 4'b1111; // x=54, y=28
        pixel_data[28][55] = 4'b0000; // x=55, y=28
        pixel_data[28][56] = 4'b0111; // x=56, y=28
        pixel_data[28][57] = 4'b0000; // x=57, y=28
        pixel_data[28][58] = 4'b0000; // x=58, y=28
        pixel_data[28][59] = 4'b0111; // x=59, y=28
        pixel_data[28][60] = 4'b1000; // x=60, y=28
        pixel_data[28][61] = 4'b1101; // x=61, y=28
        pixel_data[28][62] = 4'b0001; // x=62, y=28
        pixel_data[28][63] = 4'b1101; // x=63, y=28
        pixel_data[28][64] = 4'b0001; // x=64, y=28
        pixel_data[28][65] = 4'b1101; // x=65, y=28
        pixel_data[28][66] = 4'b0010; // x=66, y=28
        pixel_data[28][67] = 4'b0111; // x=67, y=28
        pixel_data[28][68] = 4'b0111; // x=68, y=28
        pixel_data[28][69] = 4'b0111; // x=69, y=28
        pixel_data[28][70] = 4'b0111; // x=70, y=28
        pixel_data[28][71] = 4'b0111; // x=71, y=28
        pixel_data[28][72] = 4'b0111; // x=72, y=28
        pixel_data[28][73] = 4'b0111; // x=73, y=28
        pixel_data[28][74] = 4'b0111; // x=74, y=28
        pixel_data[28][75] = 4'b1001; // x=75, y=28
        pixel_data[28][76] = 4'b1011; // x=76, y=28
        pixel_data[28][77] = 4'b0001; // x=77, y=28
        pixel_data[28][78] = 4'b0001; // x=78, y=28
        pixel_data[28][79] = 4'b0001; // x=79, y=28
        pixel_data[28][80] = 4'b1101; // x=80, y=28
        pixel_data[28][81] = 4'b0011; // x=81, y=28
        pixel_data[28][82] = 4'b1110; // x=82, y=28
        pixel_data[28][83] = 4'b0111; // x=83, y=28
        pixel_data[28][84] = 4'b0000; // x=84, y=28
        pixel_data[28][85] = 4'b0000; // x=85, y=28
        pixel_data[28][86] = 4'b0111; // x=86, y=28
        pixel_data[28][87] = 4'b0110; // x=87, y=28
        pixel_data[28][88] = 4'b1011; // x=88, y=28
        pixel_data[28][89] = 4'b1101; // x=89, y=28
        pixel_data[28][90] = 4'b1101; // x=90, y=28
        pixel_data[28][91] = 4'b1101; // x=91, y=28
        pixel_data[28][92] = 4'b1101; // x=92, y=28
        pixel_data[28][93] = 4'b0001; // x=93, y=28
        pixel_data[28][94] = 4'b1011; // x=94, y=28
        pixel_data[28][95] = 4'b0010; // x=95, y=28
        pixel_data[28][96] = 4'b1110; // x=96, y=28
        pixel_data[28][97] = 4'b0111; // x=97, y=28
        pixel_data[28][98] = 4'b0111; // x=98, y=28
        pixel_data[28][99] = 4'b0111; // x=99, y=28
        pixel_data[28][100] = 4'b0000; // x=100, y=28
        pixel_data[28][101] = 4'b0000; // x=101, y=28
        pixel_data[28][102] = 4'b0111; // x=102, y=28
        pixel_data[28][103] = 4'b0111; // x=103, y=28
        pixel_data[28][104] = 4'b0100; // x=104, y=28
        pixel_data[28][105] = 4'b0001; // x=105, y=28
        pixel_data[28][106] = 4'b0001; // x=106, y=28
        pixel_data[28][107] = 4'b0001; // x=107, y=28
        pixel_data[28][108] = 4'b0001; // x=108, y=28
        pixel_data[28][109] = 4'b1101; // x=109, y=28
        pixel_data[28][110] = 4'b1010; // x=110, y=28
        pixel_data[28][111] = 4'b0111; // x=111, y=28
        pixel_data[28][112] = 4'b0111; // x=112, y=28
        pixel_data[28][113] = 4'b0111; // x=113, y=28
        pixel_data[28][114] = 4'b0000; // x=114, y=28
        pixel_data[28][115] = 4'b0000; // x=115, y=28
        pixel_data[28][116] = 4'b0000; // x=116, y=28
        pixel_data[28][117] = 4'b0111; // x=117, y=28
        pixel_data[28][118] = 4'b0111; // x=118, y=28
        pixel_data[28][119] = 4'b1001; // x=119, y=28
        pixel_data[28][120] = 4'b0001; // x=120, y=28
        pixel_data[28][121] = 4'b1101; // x=121, y=28
        pixel_data[28][122] = 4'b0001; // x=122, y=28
        pixel_data[28][123] = 4'b0001; // x=123, y=28
        pixel_data[28][124] = 4'b1101; // x=124, y=28
        pixel_data[28][125] = 4'b1001; // x=125, y=28
        pixel_data[28][126] = 4'b0111; // x=126, y=28
        pixel_data[28][127] = 4'b0000; // x=127, y=28
        pixel_data[28][128] = 4'b0111; // x=128, y=28
        pixel_data[28][129] = 4'b0111; // x=129, y=28
        pixel_data[28][130] = 4'b0111; // x=130, y=28
        pixel_data[28][131] = 4'b0111; // x=131, y=28
        pixel_data[28][132] = 4'b0111; // x=132, y=28
        pixel_data[28][133] = 4'b0111; // x=133, y=28
        pixel_data[28][134] = 4'b0111; // x=134, y=28
        pixel_data[28][135] = 4'b0111; // x=135, y=28
        pixel_data[28][136] = 4'b0111; // x=136, y=28
        pixel_data[28][137] = 4'b0111; // x=137, y=28
        pixel_data[28][138] = 4'b0111; // x=138, y=28
        pixel_data[28][139] = 4'b0111; // x=139, y=28
        pixel_data[28][140] = 4'b0111; // x=140, y=28
        pixel_data[28][141] = 4'b0111; // x=141, y=28
        pixel_data[28][142] = 4'b0111; // x=142, y=28
        pixel_data[28][143] = 4'b1110; // x=143, y=28
        pixel_data[28][144] = 4'b1010; // x=144, y=28
        pixel_data[28][145] = 4'b0101; // x=145, y=28
        pixel_data[28][146] = 4'b0010; // x=146, y=28
        pixel_data[28][147] = 4'b0110; // x=147, y=28
        pixel_data[28][148] = 4'b0111; // x=148, y=28
        pixel_data[28][149] = 4'b0111; // x=149, y=28
        pixel_data[28][150] = 4'b0111; // x=150, y=28
        pixel_data[28][151] = 4'b0111; // x=151, y=28
        pixel_data[28][152] = 4'b0111; // x=152, y=28
        pixel_data[28][153] = 4'b0111; // x=153, y=28
        pixel_data[28][154] = 4'b0111; // x=154, y=28
        pixel_data[28][155] = 4'b0111; // x=155, y=28
        pixel_data[28][156] = 4'b0111; // x=156, y=28
        pixel_data[28][157] = 4'b0111; // x=157, y=28
        pixel_data[28][158] = 4'b0111; // x=158, y=28
        pixel_data[28][159] = 4'b0111; // x=159, y=28
        pixel_data[28][160] = 4'b0111; // x=160, y=28
        pixel_data[28][161] = 4'b0111; // x=161, y=28
        pixel_data[28][162] = 4'b0111; // x=162, y=28
        pixel_data[28][163] = 4'b0111; // x=163, y=28
        pixel_data[28][164] = 4'b0111; // x=164, y=28
        pixel_data[28][165] = 4'b0111; // x=165, y=28
        pixel_data[28][166] = 4'b0111; // x=166, y=28
        pixel_data[28][167] = 4'b0111; // x=167, y=28
        pixel_data[28][168] = 4'b0111; // x=168, y=28
        pixel_data[28][169] = 4'b0111; // x=169, y=28
        pixel_data[28][170] = 4'b0111; // x=170, y=28
        pixel_data[28][171] = 4'b0111; // x=171, y=28
        pixel_data[28][172] = 4'b0111; // x=172, y=28
        pixel_data[28][173] = 4'b0111; // x=173, y=28
        pixel_data[28][174] = 4'b0111; // x=174, y=28
        pixel_data[28][175] = 4'b0111; // x=175, y=28
        pixel_data[28][176] = 4'b0111; // x=176, y=28
        pixel_data[28][177] = 4'b0111; // x=177, y=28
        pixel_data[28][178] = 4'b0111; // x=178, y=28
        pixel_data[28][179] = 4'b0111; // x=179, y=28
        pixel_data[29][0] = 4'b0111; // x=0, y=29
        pixel_data[29][1] = 4'b0111; // x=1, y=29
        pixel_data[29][2] = 4'b0111; // x=2, y=29
        pixel_data[29][3] = 4'b0111; // x=3, y=29
        pixel_data[29][4] = 4'b0111; // x=4, y=29
        pixel_data[29][5] = 4'b0111; // x=5, y=29
        pixel_data[29][6] = 4'b0111; // x=6, y=29
        pixel_data[29][7] = 4'b0111; // x=7, y=29
        pixel_data[29][8] = 4'b0111; // x=8, y=29
        pixel_data[29][9] = 4'b0000; // x=9, y=29
        pixel_data[29][10] = 4'b0000; // x=10, y=29
        pixel_data[29][11] = 4'b0111; // x=11, y=29
        pixel_data[29][12] = 4'b1110; // x=12, y=29
        pixel_data[29][13] = 4'b0101; // x=13, y=29
        pixel_data[29][14] = 4'b1011; // x=14, y=29
        pixel_data[29][15] = 4'b1101; // x=15, y=29
        pixel_data[29][16] = 4'b1101; // x=16, y=29
        pixel_data[29][17] = 4'b1101; // x=17, y=29
        pixel_data[29][18] = 4'b1101; // x=18, y=29
        pixel_data[29][19] = 4'b0001; // x=19, y=29
        pixel_data[29][20] = 4'b0001; // x=20, y=29
        pixel_data[29][21] = 4'b0001; // x=21, y=29
        pixel_data[29][22] = 4'b0001; // x=22, y=29
        pixel_data[29][23] = 4'b0001; // x=23, y=29
        pixel_data[29][24] = 4'b1101; // x=24, y=29
        pixel_data[29][25] = 4'b1101; // x=25, y=29
        pixel_data[29][26] = 4'b1101; // x=26, y=29
        pixel_data[29][27] = 4'b1011; // x=27, y=29
        pixel_data[29][28] = 4'b0101; // x=28, y=29
        pixel_data[29][29] = 4'b1110; // x=29, y=29
        pixel_data[29][30] = 4'b0111; // x=30, y=29
        pixel_data[29][31] = 4'b0000; // x=31, y=29
        pixel_data[29][32] = 4'b0111; // x=32, y=29
        pixel_data[29][33] = 4'b0111; // x=33, y=29
        pixel_data[29][34] = 4'b0111; // x=34, y=29
        pixel_data[29][35] = 4'b0111; // x=35, y=29
        pixel_data[29][36] = 4'b0101; // x=36, y=29
        pixel_data[29][37] = 4'b1101; // x=37, y=29
        pixel_data[29][38] = 4'b0001; // x=38, y=29
        pixel_data[29][39] = 4'b1101; // x=39, y=29
        pixel_data[29][40] = 4'b1101; // x=40, y=29
        pixel_data[29][41] = 4'b1011; // x=41, y=29
        pixel_data[29][42] = 4'b1110; // x=42, y=29
        pixel_data[29][43] = 4'b0111; // x=43, y=29
        pixel_data[29][44] = 4'b0000; // x=44, y=29
        pixel_data[29][45] = 4'b0111; // x=45, y=29
        pixel_data[29][46] = 4'b0111; // x=46, y=29
        pixel_data[29][47] = 4'b0111; // x=47, y=29
        pixel_data[29][48] = 4'b0111; // x=48, y=29
        pixel_data[29][49] = 4'b0000; // x=49, y=29
        pixel_data[29][50] = 4'b0000; // x=50, y=29
        pixel_data[29][51] = 4'b0111; // x=51, y=29
        pixel_data[29][52] = 4'b0111; // x=52, y=29
        pixel_data[29][53] = 4'b0110; // x=53, y=29
        pixel_data[29][54] = 4'b0000; // x=54, y=29
        pixel_data[29][55] = 4'b0111; // x=55, y=29
        pixel_data[29][56] = 4'b0000; // x=56, y=29
        pixel_data[29][57] = 4'b0000; // x=57, y=29
        pixel_data[29][58] = 4'b0111; // x=58, y=29
        pixel_data[29][59] = 4'b0100; // x=59, y=29
        pixel_data[29][60] = 4'b0001; // x=60, y=29
        pixel_data[29][61] = 4'b1101; // x=61, y=29
        pixel_data[29][62] = 4'b1101; // x=62, y=29
        pixel_data[29][63] = 4'b0001; // x=63, y=29
        pixel_data[29][64] = 4'b1101; // x=64, y=29
        pixel_data[29][65] = 4'b0101; // x=65, y=29
        pixel_data[29][66] = 4'b0111; // x=66, y=29
        pixel_data[29][67] = 4'b0000; // x=67, y=29
        pixel_data[29][68] = 4'b0000; // x=68, y=29
        pixel_data[29][69] = 4'b0111; // x=69, y=29
        pixel_data[29][70] = 4'b0111; // x=70, y=29
        pixel_data[29][71] = 4'b0111; // x=71, y=29
        pixel_data[29][72] = 4'b0000; // x=72, y=29
        pixel_data[29][73] = 4'b0000; // x=73, y=29
        pixel_data[29][74] = 4'b0000; // x=74, y=29
        pixel_data[29][75] = 4'b0111; // x=75, y=29
        pixel_data[29][76] = 4'b1001; // x=76, y=29
        pixel_data[29][77] = 4'b1101; // x=77, y=29
        pixel_data[29][78] = 4'b1101; // x=78, y=29
        pixel_data[29][79] = 4'b1101; // x=79, y=29
        pixel_data[29][80] = 4'b0001; // x=80, y=29
        pixel_data[29][81] = 4'b1101; // x=81, y=29
        pixel_data[29][82] = 4'b1010; // x=82, y=29
        pixel_data[29][83] = 4'b0111; // x=83, y=29
        pixel_data[29][84] = 4'b0000; // x=84, y=29
        pixel_data[29][85] = 4'b0111; // x=85, y=29
        pixel_data[29][86] = 4'b0111; // x=86, y=29
        pixel_data[29][87] = 4'b0110; // x=87, y=29
        pixel_data[29][88] = 4'b1011; // x=88, y=29
        pixel_data[29][89] = 4'b1101; // x=89, y=29
        pixel_data[29][90] = 4'b0001; // x=90, y=29
        pixel_data[29][91] = 4'b1101; // x=91, y=29
        pixel_data[29][92] = 4'b1101; // x=92, y=29
        pixel_data[29][93] = 4'b0001; // x=93, y=29
        pixel_data[29][94] = 4'b1001; // x=94, y=29
        pixel_data[29][95] = 4'b0111; // x=95, y=29
        pixel_data[29][96] = 4'b0111; // x=96, y=29
        pixel_data[29][97] = 4'b0000; // x=97, y=29
        pixel_data[29][98] = 4'b0000; // x=98, y=29
        pixel_data[29][99] = 4'b0000; // x=99, y=29
        pixel_data[29][100] = 4'b0111; // x=100, y=29
        pixel_data[29][101] = 4'b0111; // x=101, y=29
        pixel_data[29][102] = 4'b0111; // x=102, y=29
        pixel_data[29][103] = 4'b0111; // x=103, y=29
        pixel_data[29][104] = 4'b1111; // x=104, y=29
        pixel_data[29][105] = 4'b1101; // x=105, y=29
        pixel_data[29][106] = 4'b0001; // x=106, y=29
        pixel_data[29][107] = 4'b0001; // x=107, y=29
        pixel_data[29][108] = 4'b1101; // x=108, y=29
        pixel_data[29][109] = 4'b0101; // x=109, y=29
        pixel_data[29][110] = 4'b0111; // x=110, y=29
        pixel_data[29][111] = 4'b0111; // x=111, y=29
        pixel_data[29][112] = 4'b0111; // x=112, y=29
        pixel_data[29][113] = 4'b0111; // x=113, y=29
        pixel_data[29][114] = 4'b0111; // x=114, y=29
        pixel_data[29][115] = 4'b0111; // x=115, y=29
        pixel_data[29][116] = 4'b0111; // x=116, y=29
        pixel_data[29][117] = 4'b0111; // x=117, y=29
        pixel_data[29][118] = 4'b0111; // x=118, y=29
        pixel_data[29][119] = 4'b0111; // x=119, y=29
        pixel_data[29][120] = 4'b0010; // x=120, y=29
        pixel_data[29][121] = 4'b1101; // x=121, y=29
        pixel_data[29][122] = 4'b1101; // x=122, y=29
        pixel_data[29][123] = 4'b0001; // x=123, y=29
        pixel_data[29][124] = 4'b1101; // x=124, y=29
        pixel_data[29][125] = 4'b1111; // x=125, y=29
        pixel_data[29][126] = 4'b0111; // x=126, y=29
        pixel_data[29][127] = 4'b0111; // x=127, y=29
        pixel_data[29][128] = 4'b0111; // x=128, y=29
        pixel_data[29][129] = 4'b0111; // x=129, y=29
        pixel_data[29][130] = 4'b0111; // x=130, y=29
        pixel_data[29][131] = 4'b0111; // x=131, y=29
        pixel_data[29][132] = 4'b0111; // x=132, y=29
        pixel_data[29][133] = 4'b0111; // x=133, y=29
        pixel_data[29][134] = 4'b0111; // x=134, y=29
        pixel_data[29][135] = 4'b0111; // x=135, y=29
        pixel_data[29][136] = 4'b0111; // x=136, y=29
        pixel_data[29][137] = 4'b0111; // x=137, y=29
        pixel_data[29][138] = 4'b0111; // x=138, y=29
        pixel_data[29][139] = 4'b0111; // x=139, y=29
        pixel_data[29][140] = 4'b0111; // x=140, y=29
        pixel_data[29][141] = 4'b0111; // x=141, y=29
        pixel_data[29][142] = 4'b0111; // x=142, y=29
        pixel_data[29][143] = 4'b0111; // x=143, y=29
        pixel_data[29][144] = 4'b0111; // x=144, y=29
        pixel_data[29][145] = 4'b0111; // x=145, y=29
        pixel_data[29][146] = 4'b0111; // x=146, y=29
        pixel_data[29][147] = 4'b0111; // x=147, y=29
        pixel_data[29][148] = 4'b0111; // x=148, y=29
        pixel_data[29][149] = 4'b0111; // x=149, y=29
        pixel_data[29][150] = 4'b0111; // x=150, y=29
        pixel_data[29][151] = 4'b0111; // x=151, y=29
        pixel_data[29][152] = 4'b0111; // x=152, y=29
        pixel_data[29][153] = 4'b0111; // x=153, y=29
        pixel_data[29][154] = 4'b0111; // x=154, y=29
        pixel_data[29][155] = 4'b0111; // x=155, y=29
        pixel_data[29][156] = 4'b0111; // x=156, y=29
        pixel_data[29][157] = 4'b0111; // x=157, y=29
        pixel_data[29][158] = 4'b0111; // x=158, y=29
        pixel_data[29][159] = 4'b0111; // x=159, y=29
        pixel_data[29][160] = 4'b0111; // x=160, y=29
        pixel_data[29][161] = 4'b0111; // x=161, y=29
        pixel_data[29][162] = 4'b0111; // x=162, y=29
        pixel_data[29][163] = 4'b0111; // x=163, y=29
        pixel_data[29][164] = 4'b0111; // x=164, y=29
        pixel_data[29][165] = 4'b0111; // x=165, y=29
        pixel_data[29][166] = 4'b0111; // x=166, y=29
        pixel_data[29][167] = 4'b0111; // x=167, y=29
        pixel_data[29][168] = 4'b0111; // x=168, y=29
        pixel_data[29][169] = 4'b0111; // x=169, y=29
        pixel_data[29][170] = 4'b0111; // x=170, y=29
        pixel_data[29][171] = 4'b0111; // x=171, y=29
        pixel_data[29][172] = 4'b0111; // x=172, y=29
        pixel_data[29][173] = 4'b0111; // x=173, y=29
        pixel_data[29][174] = 4'b0111; // x=174, y=29
        pixel_data[29][175] = 4'b0111; // x=175, y=29
        pixel_data[29][176] = 4'b0111; // x=176, y=29
        pixel_data[29][177] = 4'b0111; // x=177, y=29
        pixel_data[29][178] = 4'b0111; // x=178, y=29
        pixel_data[29][179] = 4'b0111; // x=179, y=29
        pixel_data[30][0] = 4'b0111; // x=0, y=30
        pixel_data[30][1] = 4'b0111; // x=1, y=30
        pixel_data[30][2] = 4'b0111; // x=2, y=30
        pixel_data[30][3] = 4'b0111; // x=3, y=30
        pixel_data[30][4] = 4'b0111; // x=4, y=30
        pixel_data[30][5] = 4'b0111; // x=5, y=30
        pixel_data[30][6] = 4'b0111; // x=6, y=30
        pixel_data[30][7] = 4'b0111; // x=7, y=30
        pixel_data[30][8] = 4'b0111; // x=8, y=30
        pixel_data[30][9] = 4'b0000; // x=9, y=30
        pixel_data[30][10] = 4'b0000; // x=10, y=30
        pixel_data[30][11] = 4'b0000; // x=11, y=30
        pixel_data[30][12] = 4'b0111; // x=12, y=30
        pixel_data[30][13] = 4'b0111; // x=13, y=30
        pixel_data[30][14] = 4'b0110; // x=14, y=30
        pixel_data[30][15] = 4'b0010; // x=15, y=30
        pixel_data[30][16] = 4'b1100; // x=16, y=30
        pixel_data[30][17] = 4'b1011; // x=17, y=30
        pixel_data[30][18] = 4'b1101; // x=18, y=30
        pixel_data[30][19] = 4'b1101; // x=19, y=30
        pixel_data[30][20] = 4'b1101; // x=20, y=30
        pixel_data[30][21] = 4'b1101; // x=21, y=30
        pixel_data[30][22] = 4'b1101; // x=22, y=30
        pixel_data[30][23] = 4'b0001; // x=23, y=30
        pixel_data[30][24] = 4'b0001; // x=24, y=30
        pixel_data[30][25] = 4'b1101; // x=25, y=30
        pixel_data[30][26] = 4'b0001; // x=26, y=30
        pixel_data[30][27] = 4'b1101; // x=27, y=30
        pixel_data[30][28] = 4'b1101; // x=28, y=30
        pixel_data[30][29] = 4'b0011; // x=29, y=30
        pixel_data[30][30] = 4'b0110; // x=30, y=30
        pixel_data[30][31] = 4'b0111; // x=31, y=30
        pixel_data[30][32] = 4'b0111; // x=32, y=30
        pixel_data[30][33] = 4'b0111; // x=33, y=30
        pixel_data[30][34] = 4'b0111; // x=34, y=30
        pixel_data[30][35] = 4'b0000; // x=35, y=30
        pixel_data[30][36] = 4'b0011; // x=36, y=30
        pixel_data[30][37] = 4'b1101; // x=37, y=30
        pixel_data[30][38] = 4'b0001; // x=38, y=30
        pixel_data[30][39] = 4'b1101; // x=39, y=30
        pixel_data[30][40] = 4'b1101; // x=40, y=30
        pixel_data[30][41] = 4'b1010; // x=41, y=30
        pixel_data[30][42] = 4'b0111; // x=42, y=30
        pixel_data[30][43] = 4'b0000; // x=43, y=30
        pixel_data[30][44] = 4'b0111; // x=44, y=30
        pixel_data[30][45] = 4'b0111; // x=45, y=30
        pixel_data[30][46] = 4'b0111; // x=46, y=30
        pixel_data[30][47] = 4'b0111; // x=47, y=30
        pixel_data[30][48] = 4'b0111; // x=48, y=30
        pixel_data[30][49] = 4'b0111; // x=49, y=30
        pixel_data[30][50] = 4'b0000; // x=50, y=30
        pixel_data[30][51] = 4'b0000; // x=51, y=30
        pixel_data[30][52] = 4'b0000; // x=52, y=30
        pixel_data[30][53] = 4'b0111; // x=53, y=30
        pixel_data[30][54] = 4'b0111; // x=54, y=30
        pixel_data[30][55] = 4'b0000; // x=55, y=30
        pixel_data[30][56] = 4'b0000; // x=56, y=30
        pixel_data[30][57] = 4'b0000; // x=57, y=30
        pixel_data[30][58] = 4'b0111; // x=58, y=30
        pixel_data[30][59] = 4'b0010; // x=59, y=30
        pixel_data[30][60] = 4'b1101; // x=60, y=30
        pixel_data[30][61] = 4'b0001; // x=61, y=30
        pixel_data[30][62] = 4'b1101; // x=62, y=30
        pixel_data[30][63] = 4'b1101; // x=63, y=30
        pixel_data[30][64] = 4'b1011; // x=64, y=30
        pixel_data[30][65] = 4'b1110; // x=65, y=30
        pixel_data[30][66] = 4'b0111; // x=66, y=30
        pixel_data[30][67] = 4'b0000; // x=67, y=30
        pixel_data[30][68] = 4'b0111; // x=68, y=30
        pixel_data[30][69] = 4'b0111; // x=69, y=30
        pixel_data[30][70] = 4'b0111; // x=70, y=30
        pixel_data[30][71] = 4'b0111; // x=71, y=30
        pixel_data[30][72] = 4'b0111; // x=72, y=30
        pixel_data[30][73] = 4'b0111; // x=73, y=30
        pixel_data[30][74] = 4'b0111; // x=74, y=30
        pixel_data[30][75] = 4'b0000; // x=75, y=30
        pixel_data[30][76] = 4'b0111; // x=76, y=30
        pixel_data[30][77] = 4'b1100; // x=77, y=30
        pixel_data[30][78] = 4'b1101; // x=78, y=30
        pixel_data[30][79] = 4'b0001; // x=79, y=30
        pixel_data[30][80] = 4'b0001; // x=80, y=30
        pixel_data[30][81] = 4'b1101; // x=81, y=30
        pixel_data[30][82] = 4'b1100; // x=82, y=30
        pixel_data[30][83] = 4'b0111; // x=83, y=30
        pixel_data[30][84] = 4'b0000; // x=84, y=30
        pixel_data[30][85] = 4'b0000; // x=85, y=30
        pixel_data[30][86] = 4'b0111; // x=86, y=30
        pixel_data[30][87] = 4'b0110; // x=87, y=30
        pixel_data[30][88] = 4'b1011; // x=88, y=30
        pixel_data[30][89] = 4'b1101; // x=89, y=30
        pixel_data[30][90] = 4'b0001; // x=90, y=30
        pixel_data[30][91] = 4'b0001; // x=91, y=30
        pixel_data[30][92] = 4'b1101; // x=92, y=30
        pixel_data[30][93] = 4'b1111; // x=93, y=30
        pixel_data[30][94] = 4'b0111; // x=94, y=30
        pixel_data[30][95] = 4'b0000; // x=95, y=30
        pixel_data[30][96] = 4'b0000; // x=96, y=30
        pixel_data[30][97] = 4'b0111; // x=97, y=30
        pixel_data[30][98] = 4'b0000; // x=98, y=30
        pixel_data[30][99] = 4'b0111; // x=99, y=30
        pixel_data[30][100] = 4'b0111; // x=100, y=30
        pixel_data[30][101] = 4'b0111; // x=101, y=30
        pixel_data[30][102] = 4'b0111; // x=102, y=30
        pixel_data[30][103] = 4'b1110; // x=103, y=30
        pixel_data[30][104] = 4'b1011; // x=104, y=30
        pixel_data[30][105] = 4'b1101; // x=105, y=30
        pixel_data[30][106] = 4'b1101; // x=106, y=30
        pixel_data[30][107] = 4'b1101; // x=107, y=30
        pixel_data[30][108] = 4'b1101; // x=108, y=30
        pixel_data[30][109] = 4'b1111; // x=109, y=30
        pixel_data[30][110] = 4'b0010; // x=110, y=30
        pixel_data[30][111] = 4'b0010; // x=111, y=30
        pixel_data[30][112] = 4'b0010; // x=112, y=30
        pixel_data[30][113] = 4'b0010; // x=113, y=30
        pixel_data[30][114] = 4'b0010; // x=114, y=30
        pixel_data[30][115] = 4'b0010; // x=115, y=30
        pixel_data[30][116] = 4'b0010; // x=116, y=30
        pixel_data[30][117] = 4'b0010; // x=117, y=30
        pixel_data[30][118] = 4'b0010; // x=118, y=30
        pixel_data[30][119] = 4'b0010; // x=119, y=30
        pixel_data[30][120] = 4'b1111; // x=120, y=30
        pixel_data[30][121] = 4'b0001; // x=121, y=30
        pixel_data[30][122] = 4'b1101; // x=122, y=30
        pixel_data[30][123] = 4'b1101; // x=123, y=30
        pixel_data[30][124] = 4'b1101; // x=124, y=30
        pixel_data[30][125] = 4'b0011; // x=125, y=30
        pixel_data[30][126] = 4'b0000; // x=126, y=30
        pixel_data[30][127] = 4'b0111; // x=127, y=30
        pixel_data[30][128] = 4'b0111; // x=128, y=30
        pixel_data[30][129] = 4'b0111; // x=129, y=30
        pixel_data[30][130] = 4'b0111; // x=130, y=30
        pixel_data[30][131] = 4'b0111; // x=131, y=30
        pixel_data[30][132] = 4'b0111; // x=132, y=30
        pixel_data[30][133] = 4'b0111; // x=133, y=30
        pixel_data[30][134] = 4'b0111; // x=134, y=30
        pixel_data[30][135] = 4'b0111; // x=135, y=30
        pixel_data[30][136] = 4'b0111; // x=136, y=30
        pixel_data[30][137] = 4'b0111; // x=137, y=30
        pixel_data[30][138] = 4'b0111; // x=138, y=30
        pixel_data[30][139] = 4'b0111; // x=139, y=30
        pixel_data[30][140] = 4'b0111; // x=140, y=30
        pixel_data[30][141] = 4'b0111; // x=141, y=30
        pixel_data[30][142] = 4'b0111; // x=142, y=30
        pixel_data[30][143] = 4'b0111; // x=143, y=30
        pixel_data[30][144] = 4'b0000; // x=144, y=30
        pixel_data[30][145] = 4'b0000; // x=145, y=30
        pixel_data[30][146] = 4'b0000; // x=146, y=30
        pixel_data[30][147] = 4'b0000; // x=147, y=30
        pixel_data[30][148] = 4'b0000; // x=148, y=30
        pixel_data[30][149] = 4'b0111; // x=149, y=30
        pixel_data[30][150] = 4'b0111; // x=150, y=30
        pixel_data[30][151] = 4'b0111; // x=151, y=30
        pixel_data[30][152] = 4'b0111; // x=152, y=30
        pixel_data[30][153] = 4'b0111; // x=153, y=30
        pixel_data[30][154] = 4'b0111; // x=154, y=30
        pixel_data[30][155] = 4'b0111; // x=155, y=30
        pixel_data[30][156] = 4'b0111; // x=156, y=30
        pixel_data[30][157] = 4'b0111; // x=157, y=30
        pixel_data[30][158] = 4'b0111; // x=158, y=30
        pixel_data[30][159] = 4'b0111; // x=159, y=30
        pixel_data[30][160] = 4'b0111; // x=160, y=30
        pixel_data[30][161] = 4'b0111; // x=161, y=30
        pixel_data[30][162] = 4'b0111; // x=162, y=30
        pixel_data[30][163] = 4'b0111; // x=163, y=30
        pixel_data[30][164] = 4'b0111; // x=164, y=30
        pixel_data[30][165] = 4'b0111; // x=165, y=30
        pixel_data[30][166] = 4'b0111; // x=166, y=30
        pixel_data[30][167] = 4'b0111; // x=167, y=30
        pixel_data[30][168] = 4'b0111; // x=168, y=30
        pixel_data[30][169] = 4'b0111; // x=169, y=30
        pixel_data[30][170] = 4'b0111; // x=170, y=30
        pixel_data[30][171] = 4'b0111; // x=171, y=30
        pixel_data[30][172] = 4'b0111; // x=172, y=30
        pixel_data[30][173] = 4'b0111; // x=173, y=30
        pixel_data[30][174] = 4'b0111; // x=174, y=30
        pixel_data[30][175] = 4'b0111; // x=175, y=30
        pixel_data[30][176] = 4'b0111; // x=176, y=30
        pixel_data[30][177] = 4'b0111; // x=177, y=30
        pixel_data[30][178] = 4'b0111; // x=178, y=30
        pixel_data[30][179] = 4'b0111; // x=179, y=30
        pixel_data[31][0] = 4'b0111; // x=0, y=31
        pixel_data[31][1] = 4'b0111; // x=1, y=31
        pixel_data[31][2] = 4'b0111; // x=2, y=31
        pixel_data[31][3] = 4'b0111; // x=3, y=31
        pixel_data[31][4] = 4'b0111; // x=4, y=31
        pixel_data[31][5] = 4'b0111; // x=5, y=31
        pixel_data[31][6] = 4'b0111; // x=6, y=31
        pixel_data[31][7] = 4'b0111; // x=7, y=31
        pixel_data[31][8] = 4'b0111; // x=8, y=31
        pixel_data[31][9] = 4'b0000; // x=9, y=31
        pixel_data[31][10] = 4'b0000; // x=10, y=31
        pixel_data[31][11] = 4'b0000; // x=11, y=31
        pixel_data[31][12] = 4'b0000; // x=12, y=31
        pixel_data[31][13] = 4'b0000; // x=13, y=31
        pixel_data[31][14] = 4'b0111; // x=14, y=31
        pixel_data[31][15] = 4'b0111; // x=15, y=31
        pixel_data[31][16] = 4'b0111; // x=16, y=31
        pixel_data[31][17] = 4'b1110; // x=17, y=31
        pixel_data[31][18] = 4'b0100; // x=18, y=31
        pixel_data[31][19] = 4'b1010; // x=19, y=31
        pixel_data[31][20] = 4'b1111; // x=20, y=31
        pixel_data[31][21] = 4'b1100; // x=21, y=31
        pixel_data[31][22] = 4'b1011; // x=22, y=31
        pixel_data[31][23] = 4'b1101; // x=23, y=31
        pixel_data[31][24] = 4'b1101; // x=24, y=31
        pixel_data[31][25] = 4'b0001; // x=25, y=31
        pixel_data[31][26] = 4'b1101; // x=26, y=31
        pixel_data[31][27] = 4'b1101; // x=27, y=31
        pixel_data[31][28] = 4'b0001; // x=28, y=31
        pixel_data[31][29] = 4'b1101; // x=29, y=31
        pixel_data[31][30] = 4'b0011; // x=30, y=31
        pixel_data[31][31] = 4'b1110; // x=31, y=31
        pixel_data[31][32] = 4'b0111; // x=32, y=31
        pixel_data[31][33] = 4'b0000; // x=33, y=31
        pixel_data[31][34] = 4'b0111; // x=34, y=31
        pixel_data[31][35] = 4'b1110; // x=35, y=31
        pixel_data[31][36] = 4'b0001; // x=36, y=31
        pixel_data[31][37] = 4'b1101; // x=37, y=31
        pixel_data[31][38] = 4'b0001; // x=38, y=31
        pixel_data[31][39] = 4'b1101; // x=39, y=31
        pixel_data[31][40] = 4'b1101; // x=40, y=31
        pixel_data[31][41] = 4'b0110; // x=41, y=31
        pixel_data[31][42] = 4'b0111; // x=42, y=31
        pixel_data[31][43] = 4'b0000; // x=43, y=31
        pixel_data[31][44] = 4'b0000; // x=44, y=31
        pixel_data[31][45] = 4'b0111; // x=45, y=31
        pixel_data[31][46] = 4'b0111; // x=46, y=31
        pixel_data[31][47] = 4'b0111; // x=47, y=31
        pixel_data[31][48] = 4'b0111; // x=48, y=31
        pixel_data[31][49] = 4'b0111; // x=49, y=31
        pixel_data[31][50] = 4'b0000; // x=50, y=31
        pixel_data[31][51] = 4'b0000; // x=51, y=31
        pixel_data[31][52] = 4'b0000; // x=52, y=31
        pixel_data[31][53] = 4'b0000; // x=53, y=31
        pixel_data[31][54] = 4'b0111; // x=54, y=31
        pixel_data[31][55] = 4'b0111; // x=55, y=31
        pixel_data[31][56] = 4'b0111; // x=56, y=31
        pixel_data[31][57] = 4'b0000; // x=57, y=31
        pixel_data[31][58] = 4'b0111; // x=58, y=31
        pixel_data[31][59] = 4'b1000; // x=59, y=31
        pixel_data[31][60] = 4'b1101; // x=60, y=31
        pixel_data[31][61] = 4'b0001; // x=61, y=31
        pixel_data[31][62] = 4'b0001; // x=62, y=31
        pixel_data[31][63] = 4'b1101; // x=63, y=31
        pixel_data[31][64] = 4'b1000; // x=64, y=31
        pixel_data[31][65] = 4'b0111; // x=65, y=31
        pixel_data[31][66] = 4'b0000; // x=66, y=31
        pixel_data[31][67] = 4'b0111; // x=67, y=31
        pixel_data[31][68] = 4'b0111; // x=68, y=31
        pixel_data[31][69] = 4'b0111; // x=69, y=31
        pixel_data[31][70] = 4'b0111; // x=70, y=31
        pixel_data[31][71] = 4'b0111; // x=71, y=31
        pixel_data[31][72] = 4'b0111; // x=72, y=31
        pixel_data[31][73] = 4'b0111; // x=73, y=31
        pixel_data[31][74] = 4'b0111; // x=74, y=31
        pixel_data[31][75] = 4'b0000; // x=75, y=31
        pixel_data[31][76] = 4'b0111; // x=76, y=31
        pixel_data[31][77] = 4'b0010; // x=77, y=31
        pixel_data[31][78] = 4'b1101; // x=78, y=31
        pixel_data[31][79] = 4'b0001; // x=79, y=31
        pixel_data[31][80] = 4'b0001; // x=80, y=31
        pixel_data[31][81] = 4'b1101; // x=81, y=31
        pixel_data[31][82] = 4'b0011; // x=82, y=31
        pixel_data[31][83] = 4'b1110; // x=83, y=31
        pixel_data[31][84] = 4'b0111; // x=84, y=31
        pixel_data[31][85] = 4'b0000; // x=85, y=31
        pixel_data[31][86] = 4'b0111; // x=86, y=31
        pixel_data[31][87] = 4'b0110; // x=87, y=31
        pixel_data[31][88] = 4'b1011; // x=88, y=31
        pixel_data[31][89] = 4'b1101; // x=89, y=31
        pixel_data[31][90] = 4'b0001; // x=90, y=31
        pixel_data[31][91] = 4'b0001; // x=91, y=31
        pixel_data[31][92] = 4'b1101; // x=92, y=31
        pixel_data[31][93] = 4'b1010; // x=93, y=31
        pixel_data[31][94] = 4'b0111; // x=94, y=31
        pixel_data[31][95] = 4'b0000; // x=95, y=31
        pixel_data[31][96] = 4'b0111; // x=96, y=31
        pixel_data[31][97] = 4'b0000; // x=97, y=31
        pixel_data[31][98] = 4'b0111; // x=98, y=31
        pixel_data[31][99] = 4'b0111; // x=99, y=31
        pixel_data[31][100] = 4'b0111; // x=100, y=31
        pixel_data[31][101] = 4'b0111; // x=101, y=31
        pixel_data[31][102] = 4'b0111; // x=102, y=31
        pixel_data[31][103] = 4'b0110; // x=103, y=31
        pixel_data[31][104] = 4'b0001; // x=104, y=31
        pixel_data[31][105] = 4'b1101; // x=105, y=31
        pixel_data[31][106] = 4'b1101; // x=106, y=31
        pixel_data[31][107] = 4'b1101; // x=107, y=31
        pixel_data[31][108] = 4'b1101; // x=108, y=31
        pixel_data[31][109] = 4'b1101; // x=109, y=31
        pixel_data[31][110] = 4'b1101; // x=110, y=31
        pixel_data[31][111] = 4'b1101; // x=111, y=31
        pixel_data[31][112] = 4'b1101; // x=112, y=31
        pixel_data[31][113] = 4'b1101; // x=113, y=31
        pixel_data[31][114] = 4'b1101; // x=114, y=31
        pixel_data[31][115] = 4'b1101; // x=115, y=31
        pixel_data[31][116] = 4'b1101; // x=116, y=31
        pixel_data[31][117] = 4'b1101; // x=117, y=31
        pixel_data[31][118] = 4'b1101; // x=118, y=31
        pixel_data[31][119] = 4'b1101; // x=119, y=31
        pixel_data[31][120] = 4'b1101; // x=120, y=31
        pixel_data[31][121] = 4'b0001; // x=121, y=31
        pixel_data[31][122] = 4'b0001; // x=122, y=31
        pixel_data[31][123] = 4'b0001; // x=123, y=31
        pixel_data[31][124] = 4'b1101; // x=124, y=31
        pixel_data[31][125] = 4'b1011; // x=125, y=31
        pixel_data[31][126] = 4'b0000; // x=126, y=31
        pixel_data[31][127] = 4'b0111; // x=127, y=31
        pixel_data[31][128] = 4'b0111; // x=128, y=31
        pixel_data[31][129] = 4'b0111; // x=129, y=31
        pixel_data[31][130] = 4'b0111; // x=130, y=31
        pixel_data[31][131] = 4'b0111; // x=131, y=31
        pixel_data[31][132] = 4'b0111; // x=132, y=31
        pixel_data[31][133] = 4'b0111; // x=133, y=31
        pixel_data[31][134] = 4'b0111; // x=134, y=31
        pixel_data[31][135] = 4'b0111; // x=135, y=31
        pixel_data[31][136] = 4'b0111; // x=136, y=31
        pixel_data[31][137] = 4'b0111; // x=137, y=31
        pixel_data[31][138] = 4'b0111; // x=138, y=31
        pixel_data[31][139] = 4'b0111; // x=139, y=31
        pixel_data[31][140] = 4'b0111; // x=140, y=31
        pixel_data[31][141] = 4'b0111; // x=141, y=31
        pixel_data[31][142] = 4'b0111; // x=142, y=31
        pixel_data[31][143] = 4'b0111; // x=143, y=31
        pixel_data[31][144] = 4'b0111; // x=144, y=31
        pixel_data[31][145] = 4'b0111; // x=145, y=31
        pixel_data[31][146] = 4'b0111; // x=146, y=31
        pixel_data[31][147] = 4'b0000; // x=147, y=31
        pixel_data[31][148] = 4'b0111; // x=148, y=31
        pixel_data[31][149] = 4'b0111; // x=149, y=31
        pixel_data[31][150] = 4'b0111; // x=150, y=31
        pixel_data[31][151] = 4'b0111; // x=151, y=31
        pixel_data[31][152] = 4'b0111; // x=152, y=31
        pixel_data[31][153] = 4'b0111; // x=153, y=31
        pixel_data[31][154] = 4'b0111; // x=154, y=31
        pixel_data[31][155] = 4'b0111; // x=155, y=31
        pixel_data[31][156] = 4'b0111; // x=156, y=31
        pixel_data[31][157] = 4'b0111; // x=157, y=31
        pixel_data[31][158] = 4'b0111; // x=158, y=31
        pixel_data[31][159] = 4'b0111; // x=159, y=31
        pixel_data[31][160] = 4'b0111; // x=160, y=31
        pixel_data[31][161] = 4'b0111; // x=161, y=31
        pixel_data[31][162] = 4'b0111; // x=162, y=31
        pixel_data[31][163] = 4'b0111; // x=163, y=31
        pixel_data[31][164] = 4'b0111; // x=164, y=31
        pixel_data[31][165] = 4'b0111; // x=165, y=31
        pixel_data[31][166] = 4'b0111; // x=166, y=31
        pixel_data[31][167] = 4'b0111; // x=167, y=31
        pixel_data[31][168] = 4'b0111; // x=168, y=31
        pixel_data[31][169] = 4'b0111; // x=169, y=31
        pixel_data[31][170] = 4'b0111; // x=170, y=31
        pixel_data[31][171] = 4'b0111; // x=171, y=31
        pixel_data[31][172] = 4'b0111; // x=172, y=31
        pixel_data[31][173] = 4'b0111; // x=173, y=31
        pixel_data[31][174] = 4'b0111; // x=174, y=31
        pixel_data[31][175] = 4'b0111; // x=175, y=31
        pixel_data[31][176] = 4'b0111; // x=176, y=31
        pixel_data[31][177] = 4'b0111; // x=177, y=31
        pixel_data[31][178] = 4'b0111; // x=178, y=31
        pixel_data[31][179] = 4'b0111; // x=179, y=31
        pixel_data[32][0] = 4'b0111; // x=0, y=32
        pixel_data[32][1] = 4'b0111; // x=1, y=32
        pixel_data[32][2] = 4'b0111; // x=2, y=32
        pixel_data[32][3] = 4'b0111; // x=3, y=32
        pixel_data[32][4] = 4'b0111; // x=4, y=32
        pixel_data[32][5] = 4'b0111; // x=5, y=32
        pixel_data[32][6] = 4'b0111; // x=6, y=32
        pixel_data[32][7] = 4'b0111; // x=7, y=32
        pixel_data[32][8] = 4'b0111; // x=8, y=32
        pixel_data[32][9] = 4'b0111; // x=9, y=32
        pixel_data[32][10] = 4'b0000; // x=10, y=32
        pixel_data[32][11] = 4'b0000; // x=11, y=32
        pixel_data[32][12] = 4'b0111; // x=12, y=32
        pixel_data[32][13] = 4'b0111; // x=13, y=32
        pixel_data[32][14] = 4'b0111; // x=14, y=32
        pixel_data[32][15] = 4'b0000; // x=15, y=32
        pixel_data[32][16] = 4'b0111; // x=16, y=32
        pixel_data[32][17] = 4'b0111; // x=17, y=32
        pixel_data[32][18] = 4'b0111; // x=18, y=32
        pixel_data[32][19] = 4'b0111; // x=19, y=32
        pixel_data[32][20] = 4'b0111; // x=20, y=32
        pixel_data[32][21] = 4'b0111; // x=21, y=32
        pixel_data[32][22] = 4'b0110; // x=22, y=32
        pixel_data[32][23] = 4'b1010; // x=23, y=32
        pixel_data[32][24] = 4'b0011; // x=24, y=32
        pixel_data[32][25] = 4'b1101; // x=25, y=32
        pixel_data[32][26] = 4'b0001; // x=26, y=32
        pixel_data[32][27] = 4'b1101; // x=27, y=32
        pixel_data[32][28] = 4'b1101; // x=28, y=32
        pixel_data[32][29] = 4'b0001; // x=29, y=32
        pixel_data[32][30] = 4'b1101; // x=30, y=32
        pixel_data[32][31] = 4'b0101; // x=31, y=32
        pixel_data[32][32] = 4'b0111; // x=32, y=32
        pixel_data[32][33] = 4'b0000; // x=33, y=32
        pixel_data[32][34] = 4'b0111; // x=34, y=32
        pixel_data[32][35] = 4'b0110; // x=35, y=32
        pixel_data[32][36] = 4'b0001; // x=36, y=32
        pixel_data[32][37] = 4'b1101; // x=37, y=32
        pixel_data[32][38] = 4'b1101; // x=38, y=32
        pixel_data[32][39] = 4'b1101; // x=39, y=32
        pixel_data[32][40] = 4'b0001; // x=40, y=32
        pixel_data[32][41] = 4'b1110; // x=41, y=32
        pixel_data[32][42] = 4'b0111; // x=42, y=32
        pixel_data[32][43] = 4'b0000; // x=43, y=32
        pixel_data[32][44] = 4'b0111; // x=44, y=32
        pixel_data[32][45] = 4'b0111; // x=45, y=32
        pixel_data[32][46] = 4'b0111; // x=46, y=32
        pixel_data[32][47] = 4'b0111; // x=47, y=32
        pixel_data[32][48] = 4'b0111; // x=48, y=32
        pixel_data[32][49] = 4'b0111; // x=49, y=32
        pixel_data[32][50] = 4'b0111; // x=50, y=32
        pixel_data[32][51] = 4'b0111; // x=51, y=32
        pixel_data[32][52] = 4'b0111; // x=52, y=32
        pixel_data[32][53] = 4'b0111; // x=53, y=32
        pixel_data[32][54] = 4'b0111; // x=54, y=32
        pixel_data[32][55] = 4'b0111; // x=55, y=32
        pixel_data[32][56] = 4'b0111; // x=56, y=32
        pixel_data[32][57] = 4'b0111; // x=57, y=32
        pixel_data[32][58] = 4'b0111; // x=58, y=32
        pixel_data[32][59] = 4'b1100; // x=59, y=32
        pixel_data[32][60] = 4'b1101; // x=60, y=32
        pixel_data[32][61] = 4'b0001; // x=61, y=32
        pixel_data[32][62] = 4'b0001; // x=62, y=32
        pixel_data[32][63] = 4'b1101; // x=63, y=32
        pixel_data[32][64] = 4'b1111; // x=64, y=32
        pixel_data[32][65] = 4'b0111; // x=65, y=32
        pixel_data[32][66] = 4'b0000; // x=66, y=32
        pixel_data[32][67] = 4'b0111; // x=67, y=32
        pixel_data[32][68] = 4'b0111; // x=68, y=32
        pixel_data[32][69] = 4'b0111; // x=69, y=32
        pixel_data[32][70] = 4'b0111; // x=70, y=32
        pixel_data[32][71] = 4'b0111; // x=71, y=32
        pixel_data[32][72] = 4'b0111; // x=72, y=32
        pixel_data[32][73] = 4'b0111; // x=73, y=32
        pixel_data[32][74] = 4'b0111; // x=74, y=32
        pixel_data[32][75] = 4'b0000; // x=75, y=32
        pixel_data[32][76] = 4'b0111; // x=76, y=32
        pixel_data[32][77] = 4'b1010; // x=77, y=32
        pixel_data[32][78] = 4'b1101; // x=78, y=32
        pixel_data[32][79] = 4'b0001; // x=79, y=32
        pixel_data[32][80] = 4'b0001; // x=80, y=32
        pixel_data[32][81] = 4'b1101; // x=81, y=32
        pixel_data[32][82] = 4'b1011; // x=82, y=32
        pixel_data[32][83] = 4'b1110; // x=83, y=32
        pixel_data[32][84] = 4'b0111; // x=84, y=32
        pixel_data[32][85] = 4'b0000; // x=85, y=32
        pixel_data[32][86] = 4'b0111; // x=86, y=32
        pixel_data[32][87] = 4'b0110; // x=87, y=32
        pixel_data[32][88] = 4'b1011; // x=88, y=32
        pixel_data[32][89] = 4'b1101; // x=89, y=32
        pixel_data[32][90] = 4'b0001; // x=90, y=32
        pixel_data[32][91] = 4'b0001; // x=91, y=32
        pixel_data[32][92] = 4'b1101; // x=92, y=32
        pixel_data[32][93] = 4'b1001; // x=93, y=32
        pixel_data[32][94] = 4'b0111; // x=94, y=32
        pixel_data[32][95] = 4'b0000; // x=95, y=32
        pixel_data[32][96] = 4'b0111; // x=96, y=32
        pixel_data[32][97] = 4'b0111; // x=97, y=32
        pixel_data[32][98] = 4'b0111; // x=98, y=32
        pixel_data[32][99] = 4'b0111; // x=99, y=32
        pixel_data[32][100] = 4'b0111; // x=100, y=32
        pixel_data[32][101] = 4'b0000; // x=101, y=32
        pixel_data[32][102] = 4'b0111; // x=102, y=32
        pixel_data[32][103] = 4'b0100; // x=103, y=32
        pixel_data[32][104] = 4'b1101; // x=104, y=32
        pixel_data[32][105] = 4'b1101; // x=105, y=32
        pixel_data[32][106] = 4'b1101; // x=106, y=32
        pixel_data[32][107] = 4'b1101; // x=107, y=32
        pixel_data[32][108] = 4'b1101; // x=108, y=32
        pixel_data[32][109] = 4'b1101; // x=109, y=32
        pixel_data[32][110] = 4'b1101; // x=110, y=32
        pixel_data[32][111] = 4'b1101; // x=111, y=32
        pixel_data[32][112] = 4'b1101; // x=112, y=32
        pixel_data[32][113] = 4'b1101; // x=113, y=32
        pixel_data[32][114] = 4'b1101; // x=114, y=32
        pixel_data[32][115] = 4'b1101; // x=115, y=32
        pixel_data[32][116] = 4'b1101; // x=116, y=32
        pixel_data[32][117] = 4'b1101; // x=117, y=32
        pixel_data[32][118] = 4'b1101; // x=118, y=32
        pixel_data[32][119] = 4'b1101; // x=119, y=32
        pixel_data[32][120] = 4'b1101; // x=120, y=32
        pixel_data[32][121] = 4'b1101; // x=121, y=32
        pixel_data[32][122] = 4'b1101; // x=122, y=32
        pixel_data[32][123] = 4'b1101; // x=123, y=32
        pixel_data[32][124] = 4'b1101; // x=124, y=32
        pixel_data[32][125] = 4'b0001; // x=125, y=32
        pixel_data[32][126] = 4'b0000; // x=126, y=32
        pixel_data[32][127] = 4'b0111; // x=127, y=32
        pixel_data[32][128] = 4'b0111; // x=128, y=32
        pixel_data[32][129] = 4'b0111; // x=129, y=32
        pixel_data[32][130] = 4'b0111; // x=130, y=32
        pixel_data[32][131] = 4'b0111; // x=131, y=32
        pixel_data[32][132] = 4'b0111; // x=132, y=32
        pixel_data[32][133] = 4'b0111; // x=133, y=32
        pixel_data[32][134] = 4'b0111; // x=134, y=32
        pixel_data[32][135] = 4'b0111; // x=135, y=32
        pixel_data[32][136] = 4'b0111; // x=136, y=32
        pixel_data[32][137] = 4'b0111; // x=137, y=32
        pixel_data[32][138] = 4'b0111; // x=138, y=32
        pixel_data[32][139] = 4'b0111; // x=139, y=32
        pixel_data[32][140] = 4'b0111; // x=140, y=32
        pixel_data[32][141] = 4'b0111; // x=141, y=32
        pixel_data[32][142] = 4'b0111; // x=142, y=32
        pixel_data[32][143] = 4'b0111; // x=143, y=32
        pixel_data[32][144] = 4'b0111; // x=144, y=32
        pixel_data[32][145] = 4'b0111; // x=145, y=32
        pixel_data[32][146] = 4'b0111; // x=146, y=32
        pixel_data[32][147] = 4'b0111; // x=147, y=32
        pixel_data[32][148] = 4'b0111; // x=148, y=32
        pixel_data[32][149] = 4'b0111; // x=149, y=32
        pixel_data[32][150] = 4'b0111; // x=150, y=32
        pixel_data[32][151] = 4'b0111; // x=151, y=32
        pixel_data[32][152] = 4'b0111; // x=152, y=32
        pixel_data[32][153] = 4'b0111; // x=153, y=32
        pixel_data[32][154] = 4'b0111; // x=154, y=32
        pixel_data[32][155] = 4'b0111; // x=155, y=32
        pixel_data[32][156] = 4'b0111; // x=156, y=32
        pixel_data[32][157] = 4'b0111; // x=157, y=32
        pixel_data[32][158] = 4'b0111; // x=158, y=32
        pixel_data[32][159] = 4'b0111; // x=159, y=32
        pixel_data[32][160] = 4'b0111; // x=160, y=32
        pixel_data[32][161] = 4'b0111; // x=161, y=32
        pixel_data[32][162] = 4'b0111; // x=162, y=32
        pixel_data[32][163] = 4'b0111; // x=163, y=32
        pixel_data[32][164] = 4'b0111; // x=164, y=32
        pixel_data[32][165] = 4'b0111; // x=165, y=32
        pixel_data[32][166] = 4'b0111; // x=166, y=32
        pixel_data[32][167] = 4'b0111; // x=167, y=32
        pixel_data[32][168] = 4'b0111; // x=168, y=32
        pixel_data[32][169] = 4'b0111; // x=169, y=32
        pixel_data[32][170] = 4'b0111; // x=170, y=32
        pixel_data[32][171] = 4'b0111; // x=171, y=32
        pixel_data[32][172] = 4'b0111; // x=172, y=32
        pixel_data[32][173] = 4'b0111; // x=173, y=32
        pixel_data[32][174] = 4'b0111; // x=174, y=32
        pixel_data[32][175] = 4'b0111; // x=175, y=32
        pixel_data[32][176] = 4'b0111; // x=176, y=32
        pixel_data[32][177] = 4'b0111; // x=177, y=32
        pixel_data[32][178] = 4'b0111; // x=178, y=32
        pixel_data[32][179] = 4'b0111; // x=179, y=32
        pixel_data[33][0] = 4'b0111; // x=0, y=33
        pixel_data[33][1] = 4'b0111; // x=1, y=33
        pixel_data[33][2] = 4'b0111; // x=2, y=33
        pixel_data[33][3] = 4'b0111; // x=3, y=33
        pixel_data[33][4] = 4'b0111; // x=4, y=33
        pixel_data[33][5] = 4'b0111; // x=5, y=33
        pixel_data[33][6] = 4'b0111; // x=6, y=33
        pixel_data[33][7] = 4'b0111; // x=7, y=33
        pixel_data[33][8] = 4'b0111; // x=8, y=33
        pixel_data[33][9] = 4'b0000; // x=9, y=33
        pixel_data[33][10] = 4'b0000; // x=10, y=33
        pixel_data[33][11] = 4'b0111; // x=11, y=33
        pixel_data[33][12] = 4'b0000; // x=12, y=33
        pixel_data[33][13] = 4'b0111; // x=13, y=33
        pixel_data[33][14] = 4'b0111; // x=14, y=33
        pixel_data[33][15] = 4'b0111; // x=15, y=33
        pixel_data[33][16] = 4'b0111; // x=16, y=33
        pixel_data[33][17] = 4'b0111; // x=17, y=33
        pixel_data[33][18] = 4'b0000; // x=18, y=33
        pixel_data[33][19] = 4'b0000; // x=19, y=33
        pixel_data[33][20] = 4'b0000; // x=20, y=33
        pixel_data[33][21] = 4'b0000; // x=21, y=33
        pixel_data[33][22] = 4'b0111; // x=22, y=33
        pixel_data[33][23] = 4'b0111; // x=23, y=33
        pixel_data[33][24] = 4'b0000; // x=24, y=33
        pixel_data[33][25] = 4'b0101; // x=25, y=33
        pixel_data[33][26] = 4'b1101; // x=26, y=33
        pixel_data[33][27] = 4'b1101; // x=27, y=33
        pixel_data[33][28] = 4'b1101; // x=28, y=33
        pixel_data[33][29] = 4'b0001; // x=29, y=33
        pixel_data[33][30] = 4'b1101; // x=30, y=33
        pixel_data[33][31] = 4'b1100; // x=31, y=33
        pixel_data[33][32] = 4'b0000; // x=32, y=33
        pixel_data[33][33] = 4'b0111; // x=33, y=33
        pixel_data[33][34] = 4'b0111; // x=34, y=33
        pixel_data[33][35] = 4'b1110; // x=35, y=33
        pixel_data[33][36] = 4'b0001; // x=36, y=33
        pixel_data[33][37] = 4'b1101; // x=37, y=33
        pixel_data[33][38] = 4'b1101; // x=38, y=33
        pixel_data[33][39] = 4'b1101; // x=39, y=33
        pixel_data[33][40] = 4'b1101; // x=40, y=33
        pixel_data[33][41] = 4'b0110; // x=41, y=33
        pixel_data[33][42] = 4'b0111; // x=42, y=33
        pixel_data[33][43] = 4'b0000; // x=43, y=33
        pixel_data[33][44] = 4'b0111; // x=44, y=33
        pixel_data[33][45] = 4'b0111; // x=45, y=33
        pixel_data[33][46] = 4'b0111; // x=46, y=33
        pixel_data[33][47] = 4'b0111; // x=47, y=33
        pixel_data[33][48] = 4'b0111; // x=48, y=33
        pixel_data[33][49] = 4'b0111; // x=49, y=33
        pixel_data[33][50] = 4'b0111; // x=50, y=33
        pixel_data[33][51] = 4'b0111; // x=51, y=33
        pixel_data[33][52] = 4'b0111; // x=52, y=33
        pixel_data[33][53] = 4'b0111; // x=53, y=33
        pixel_data[33][54] = 4'b0111; // x=54, y=33
        pixel_data[33][55] = 4'b0111; // x=55, y=33
        pixel_data[33][56] = 4'b0111; // x=56, y=33
        pixel_data[33][57] = 4'b0111; // x=57, y=33
        pixel_data[33][58] = 4'b0111; // x=58, y=33
        pixel_data[33][59] = 4'b1000; // x=59, y=33
        pixel_data[33][60] = 4'b1101; // x=60, y=33
        pixel_data[33][61] = 4'b1101; // x=61, y=33
        pixel_data[33][62] = 4'b0001; // x=62, y=33
        pixel_data[33][63] = 4'b1101; // x=63, y=33
        pixel_data[33][64] = 4'b1100; // x=64, y=33
        pixel_data[33][65] = 4'b0111; // x=65, y=33
        pixel_data[33][66] = 4'b0000; // x=66, y=33
        pixel_data[33][67] = 4'b0111; // x=67, y=33
        pixel_data[33][68] = 4'b0111; // x=68, y=33
        pixel_data[33][69] = 4'b0111; // x=69, y=33
        pixel_data[33][70] = 4'b0111; // x=70, y=33
        pixel_data[33][71] = 4'b0111; // x=71, y=33
        pixel_data[33][72] = 4'b0111; // x=72, y=33
        pixel_data[33][73] = 4'b0111; // x=73, y=33
        pixel_data[33][74] = 4'b0111; // x=74, y=33
        pixel_data[33][75] = 4'b0000; // x=75, y=33
        pixel_data[33][76] = 4'b0111; // x=76, y=33
        pixel_data[33][77] = 4'b0101; // x=77, y=33
        pixel_data[33][78] = 4'b1101; // x=78, y=33
        pixel_data[33][79] = 4'b0001; // x=79, y=33
        pixel_data[33][80] = 4'b0001; // x=80, y=33
        pixel_data[33][81] = 4'b1101; // x=81, y=33
        pixel_data[33][82] = 4'b0011; // x=82, y=33
        pixel_data[33][83] = 4'b0000; // x=83, y=33
        pixel_data[33][84] = 4'b0111; // x=84, y=33
        pixel_data[33][85] = 4'b0000; // x=85, y=33
        pixel_data[33][86] = 4'b0111; // x=86, y=33
        pixel_data[33][87] = 4'b0110; // x=87, y=33
        pixel_data[33][88] = 4'b1011; // x=88, y=33
        pixel_data[33][89] = 4'b1101; // x=89, y=33
        pixel_data[33][90] = 4'b0001; // x=90, y=33
        pixel_data[33][91] = 4'b0001; // x=91, y=33
        pixel_data[33][92] = 4'b1101; // x=92, y=33
        pixel_data[33][93] = 4'b1001; // x=93, y=33
        pixel_data[33][94] = 4'b0111; // x=94, y=33
        pixel_data[33][95] = 4'b0000; // x=95, y=33
        pixel_data[33][96] = 4'b0111; // x=96, y=33
        pixel_data[33][97] = 4'b0111; // x=97, y=33
        pixel_data[33][98] = 4'b0111; // x=98, y=33
        pixel_data[33][99] = 4'b0111; // x=99, y=33
        pixel_data[33][100] = 4'b0111; // x=100, y=33
        pixel_data[33][101] = 4'b0111; // x=101, y=33
        pixel_data[33][102] = 4'b0111; // x=102, y=33
        pixel_data[33][103] = 4'b0110; // x=103, y=33
        pixel_data[33][104] = 4'b0001; // x=104, y=33
        pixel_data[33][105] = 4'b1101; // x=105, y=33
        pixel_data[33][106] = 4'b1101; // x=106, y=33
        pixel_data[33][107] = 4'b1101; // x=107, y=33
        pixel_data[33][108] = 4'b1101; // x=108, y=33
        pixel_data[33][109] = 4'b0010; // x=109, y=33
        pixel_data[33][110] = 4'b1010; // x=110, y=33
        pixel_data[33][111] = 4'b1010; // x=111, y=33
        pixel_data[33][112] = 4'b1010; // x=112, y=33
        pixel_data[33][113] = 4'b1010; // x=113, y=33
        pixel_data[33][114] = 4'b1010; // x=114, y=33
        pixel_data[33][115] = 4'b1010; // x=115, y=33
        pixel_data[33][116] = 4'b1010; // x=116, y=33
        pixel_data[33][117] = 4'b1010; // x=117, y=33
        pixel_data[33][118] = 4'b1010; // x=118, y=33
        pixel_data[33][119] = 4'b1010; // x=119, y=33
        pixel_data[33][120] = 4'b1010; // x=120, y=33
        pixel_data[33][121] = 4'b1010; // x=121, y=33
        pixel_data[33][122] = 4'b1010; // x=122, y=33
        pixel_data[33][123] = 4'b1010; // x=123, y=33
        pixel_data[33][124] = 4'b1010; // x=124, y=33
        pixel_data[33][125] = 4'b1010; // x=125, y=33
        pixel_data[33][126] = 4'b0000; // x=126, y=33
        pixel_data[33][127] = 4'b0111; // x=127, y=33
        pixel_data[33][128] = 4'b0111; // x=128, y=33
        pixel_data[33][129] = 4'b0111; // x=129, y=33
        pixel_data[33][130] = 4'b0111; // x=130, y=33
        pixel_data[33][131] = 4'b0111; // x=131, y=33
        pixel_data[33][132] = 4'b0111; // x=132, y=33
        pixel_data[33][133] = 4'b0111; // x=133, y=33
        pixel_data[33][134] = 4'b0111; // x=134, y=33
        pixel_data[33][135] = 4'b0111; // x=135, y=33
        pixel_data[33][136] = 4'b0111; // x=136, y=33
        pixel_data[33][137] = 4'b0111; // x=137, y=33
        pixel_data[33][138] = 4'b0111; // x=138, y=33
        pixel_data[33][139] = 4'b0111; // x=139, y=33
        pixel_data[33][140] = 4'b0111; // x=140, y=33
        pixel_data[33][141] = 4'b0111; // x=141, y=33
        pixel_data[33][142] = 4'b0111; // x=142, y=33
        pixel_data[33][143] = 4'b0111; // x=143, y=33
        pixel_data[33][144] = 4'b0111; // x=144, y=33
        pixel_data[33][145] = 4'b0111; // x=145, y=33
        pixel_data[33][146] = 4'b0111; // x=146, y=33
        pixel_data[33][147] = 4'b0111; // x=147, y=33
        pixel_data[33][148] = 4'b0111; // x=148, y=33
        pixel_data[33][149] = 4'b0111; // x=149, y=33
        pixel_data[33][150] = 4'b0111; // x=150, y=33
        pixel_data[33][151] = 4'b0111; // x=151, y=33
        pixel_data[33][152] = 4'b0111; // x=152, y=33
        pixel_data[33][153] = 4'b0111; // x=153, y=33
        pixel_data[33][154] = 4'b0111; // x=154, y=33
        pixel_data[33][155] = 4'b0111; // x=155, y=33
        pixel_data[33][156] = 4'b0111; // x=156, y=33
        pixel_data[33][157] = 4'b0111; // x=157, y=33
        pixel_data[33][158] = 4'b0111; // x=158, y=33
        pixel_data[33][159] = 4'b0111; // x=159, y=33
        pixel_data[33][160] = 4'b0111; // x=160, y=33
        pixel_data[33][161] = 4'b0111; // x=161, y=33
        pixel_data[33][162] = 4'b0111; // x=162, y=33
        pixel_data[33][163] = 4'b0111; // x=163, y=33
        pixel_data[33][164] = 4'b0111; // x=164, y=33
        pixel_data[33][165] = 4'b0111; // x=165, y=33
        pixel_data[33][166] = 4'b0111; // x=166, y=33
        pixel_data[33][167] = 4'b0111; // x=167, y=33
        pixel_data[33][168] = 4'b0111; // x=168, y=33
        pixel_data[33][169] = 4'b0111; // x=169, y=33
        pixel_data[33][170] = 4'b0111; // x=170, y=33
        pixel_data[33][171] = 4'b0111; // x=171, y=33
        pixel_data[33][172] = 4'b0111; // x=172, y=33
        pixel_data[33][173] = 4'b0111; // x=173, y=33
        pixel_data[33][174] = 4'b0111; // x=174, y=33
        pixel_data[33][175] = 4'b0111; // x=175, y=33
        pixel_data[33][176] = 4'b0111; // x=176, y=33
        pixel_data[33][177] = 4'b0111; // x=177, y=33
        pixel_data[33][178] = 4'b0111; // x=178, y=33
        pixel_data[33][179] = 4'b0111; // x=179, y=33
        pixel_data[34][0] = 4'b0111; // x=0, y=34
        pixel_data[34][1] = 4'b0111; // x=1, y=34
        pixel_data[34][2] = 4'b0111; // x=2, y=34
        pixel_data[34][3] = 4'b0111; // x=3, y=34
        pixel_data[34][4] = 4'b0111; // x=4, y=34
        pixel_data[34][5] = 4'b0111; // x=5, y=34
        pixel_data[34][6] = 4'b0111; // x=6, y=34
        pixel_data[34][7] = 4'b0111; // x=7, y=34
        pixel_data[34][8] = 4'b0111; // x=8, y=34
        pixel_data[34][9] = 4'b0111; // x=9, y=34
        pixel_data[34][10] = 4'b0111; // x=10, y=34
        pixel_data[34][11] = 4'b0101; // x=11, y=34
        pixel_data[34][12] = 4'b1100; // x=12, y=34
        pixel_data[34][13] = 4'b0000; // x=13, y=34
        pixel_data[34][14] = 4'b0111; // x=14, y=34
        pixel_data[34][15] = 4'b0000; // x=15, y=34
        pixel_data[34][16] = 4'b0111; // x=16, y=34
        pixel_data[34][17] = 4'b0111; // x=17, y=34
        pixel_data[34][18] = 4'b0000; // x=18, y=34
        pixel_data[34][19] = 4'b0111; // x=19, y=34
        pixel_data[34][20] = 4'b0111; // x=20, y=34
        pixel_data[34][21] = 4'b0111; // x=21, y=34
        pixel_data[34][22] = 4'b0000; // x=22, y=34
        pixel_data[34][23] = 4'b0000; // x=23, y=34
        pixel_data[34][24] = 4'b0111; // x=24, y=34
        pixel_data[34][25] = 4'b1110; // x=25, y=34
        pixel_data[34][26] = 4'b0011; // x=26, y=34
        pixel_data[34][27] = 4'b1101; // x=27, y=34
        pixel_data[34][28] = 4'b1101; // x=28, y=34
        pixel_data[34][29] = 4'b1101; // x=29, y=34
        pixel_data[34][30] = 4'b1101; // x=30, y=34
        pixel_data[34][31] = 4'b0011; // x=31, y=34
        pixel_data[34][32] = 4'b0000; // x=32, y=34
        pixel_data[34][33] = 4'b0111; // x=33, y=34
        pixel_data[34][34] = 4'b0111; // x=34, y=34
        pixel_data[34][35] = 4'b0000; // x=35, y=34
        pixel_data[34][36] = 4'b0011; // x=36, y=34
        pixel_data[34][37] = 4'b1101; // x=37, y=34
        pixel_data[34][38] = 4'b0001; // x=38, y=34
        pixel_data[34][39] = 4'b0001; // x=39, y=34
        pixel_data[34][40] = 4'b1101; // x=40, y=34
        pixel_data[34][41] = 4'b0010; // x=41, y=34
        pixel_data[34][42] = 4'b0111; // x=42, y=34
        pixel_data[34][43] = 4'b0000; // x=43, y=34
        pixel_data[34][44] = 4'b0111; // x=44, y=34
        pixel_data[34][45] = 4'b0111; // x=45, y=34
        pixel_data[34][46] = 4'b0111; // x=46, y=34
        pixel_data[34][47] = 4'b0111; // x=47, y=34
        pixel_data[34][48] = 4'b0111; // x=48, y=34
        pixel_data[34][49] = 4'b0111; // x=49, y=34
        pixel_data[34][50] = 4'b0111; // x=50, y=34
        pixel_data[34][51] = 4'b0111; // x=51, y=34
        pixel_data[34][52] = 4'b0000; // x=52, y=34
        pixel_data[34][53] = 4'b0111; // x=53, y=34
        pixel_data[34][54] = 4'b0111; // x=54, y=34
        pixel_data[34][55] = 4'b0111; // x=55, y=34
        pixel_data[34][56] = 4'b0111; // x=56, y=34
        pixel_data[34][57] = 4'b0000; // x=57, y=34
        pixel_data[34][58] = 4'b0111; // x=58, y=34
        pixel_data[34][59] = 4'b0010; // x=59, y=34
        pixel_data[34][60] = 4'b1101; // x=60, y=34
        pixel_data[34][61] = 4'b0001; // x=61, y=34
        pixel_data[34][62] = 4'b1101; // x=62, y=34
        pixel_data[34][63] = 4'b1101; // x=63, y=34
        pixel_data[34][64] = 4'b1011; // x=64, y=34
        pixel_data[34][65] = 4'b1110; // x=65, y=34
        pixel_data[34][66] = 4'b0111; // x=66, y=34
        pixel_data[34][67] = 4'b0000; // x=67, y=34
        pixel_data[34][68] = 4'b0111; // x=68, y=34
        pixel_data[34][69] = 4'b0111; // x=69, y=34
        pixel_data[34][70] = 4'b0111; // x=70, y=34
        pixel_data[34][71] = 4'b0111; // x=71, y=34
        pixel_data[34][72] = 4'b0111; // x=72, y=34
        pixel_data[34][73] = 4'b0111; // x=73, y=34
        pixel_data[34][74] = 4'b0111; // x=74, y=34
        pixel_data[34][75] = 4'b0000; // x=75, y=34
        pixel_data[34][76] = 4'b0111; // x=76, y=34
        pixel_data[34][77] = 4'b1100; // x=77, y=34
        pixel_data[34][78] = 4'b1101; // x=78, y=34
        pixel_data[34][79] = 4'b0001; // x=79, y=34
        pixel_data[34][80] = 4'b0001; // x=80, y=34
        pixel_data[34][81] = 4'b1101; // x=81, y=34
        pixel_data[34][82] = 4'b1000; // x=82, y=34
        pixel_data[34][83] = 4'b0111; // x=83, y=34
        pixel_data[34][84] = 4'b0000; // x=84, y=34
        pixel_data[34][85] = 4'b0111; // x=85, y=34
        pixel_data[34][86] = 4'b0111; // x=86, y=34
        pixel_data[34][87] = 4'b0110; // x=87, y=34
        pixel_data[34][88] = 4'b1011; // x=88, y=34
        pixel_data[34][89] = 4'b1101; // x=89, y=34
        pixel_data[34][90] = 4'b0001; // x=90, y=34
        pixel_data[34][91] = 4'b0001; // x=91, y=34
        pixel_data[34][92] = 4'b1101; // x=92, y=34
        pixel_data[34][93] = 4'b1001; // x=93, y=34
        pixel_data[34][94] = 4'b0111; // x=94, y=34
        pixel_data[34][95] = 4'b0000; // x=95, y=34
        pixel_data[34][96] = 4'b0111; // x=96, y=34
        pixel_data[34][97] = 4'b0111; // x=97, y=34
        pixel_data[34][98] = 4'b0111; // x=98, y=34
        pixel_data[34][99] = 4'b0111; // x=99, y=34
        pixel_data[34][100] = 4'b0111; // x=100, y=34
        pixel_data[34][101] = 4'b0111; // x=101, y=34
        pixel_data[34][102] = 4'b0111; // x=102, y=34
        pixel_data[34][103] = 4'b0000; // x=103, y=34
        pixel_data[34][104] = 4'b1011; // x=104, y=34
        pixel_data[34][105] = 4'b1101; // x=105, y=34
        pixel_data[34][106] = 4'b0001; // x=106, y=34
        pixel_data[34][107] = 4'b0001; // x=107, y=34
        pixel_data[34][108] = 4'b1101; // x=108, y=34
        pixel_data[34][109] = 4'b1010; // x=109, y=34
        pixel_data[34][110] = 4'b0111; // x=110, y=34
        pixel_data[34][111] = 4'b0111; // x=111, y=34
        pixel_data[34][112] = 4'b0111; // x=112, y=34
        pixel_data[34][113] = 4'b0111; // x=113, y=34
        pixel_data[34][114] = 4'b0111; // x=114, y=34
        pixel_data[34][115] = 4'b0111; // x=115, y=34
        pixel_data[34][116] = 4'b0111; // x=116, y=34
        pixel_data[34][117] = 4'b0111; // x=117, y=34
        pixel_data[34][118] = 4'b0111; // x=118, y=34
        pixel_data[34][119] = 4'b0111; // x=119, y=34
        pixel_data[34][120] = 4'b0111; // x=120, y=34
        pixel_data[34][121] = 4'b0111; // x=121, y=34
        pixel_data[34][122] = 4'b0111; // x=122, y=34
        pixel_data[34][123] = 4'b0111; // x=123, y=34
        pixel_data[34][124] = 4'b0111; // x=124, y=34
        pixel_data[34][125] = 4'b0111; // x=125, y=34
        pixel_data[34][126] = 4'b0111; // x=126, y=34
        pixel_data[34][127] = 4'b0111; // x=127, y=34
        pixel_data[34][128] = 4'b0111; // x=128, y=34
        pixel_data[34][129] = 4'b0111; // x=129, y=34
        pixel_data[34][130] = 4'b0111; // x=130, y=34
        pixel_data[34][131] = 4'b0111; // x=131, y=34
        pixel_data[34][132] = 4'b0111; // x=132, y=34
        pixel_data[34][133] = 4'b0111; // x=133, y=34
        pixel_data[34][134] = 4'b0111; // x=134, y=34
        pixel_data[34][135] = 4'b0111; // x=135, y=34
        pixel_data[34][136] = 4'b0111; // x=136, y=34
        pixel_data[34][137] = 4'b0111; // x=137, y=34
        pixel_data[34][138] = 4'b0111; // x=138, y=34
        pixel_data[34][139] = 4'b0111; // x=139, y=34
        pixel_data[34][140] = 4'b0111; // x=140, y=34
        pixel_data[34][141] = 4'b0111; // x=141, y=34
        pixel_data[34][142] = 4'b0111; // x=142, y=34
        pixel_data[34][143] = 4'b0111; // x=143, y=34
        pixel_data[34][144] = 4'b0000; // x=144, y=34
        pixel_data[34][145] = 4'b0000; // x=145, y=34
        pixel_data[34][146] = 4'b0000; // x=146, y=34
        pixel_data[34][147] = 4'b0000; // x=147, y=34
        pixel_data[34][148] = 4'b0111; // x=148, y=34
        pixel_data[34][149] = 4'b0111; // x=149, y=34
        pixel_data[34][150] = 4'b0111; // x=150, y=34
        pixel_data[34][151] = 4'b0111; // x=151, y=34
        pixel_data[34][152] = 4'b0111; // x=152, y=34
        pixel_data[34][153] = 4'b0111; // x=153, y=34
        pixel_data[34][154] = 4'b0111; // x=154, y=34
        pixel_data[34][155] = 4'b0111; // x=155, y=34
        pixel_data[34][156] = 4'b0111; // x=156, y=34
        pixel_data[34][157] = 4'b0111; // x=157, y=34
        pixel_data[34][158] = 4'b0111; // x=158, y=34
        pixel_data[34][159] = 4'b0111; // x=159, y=34
        pixel_data[34][160] = 4'b0111; // x=160, y=34
        pixel_data[34][161] = 4'b0111; // x=161, y=34
        pixel_data[34][162] = 4'b0111; // x=162, y=34
        pixel_data[34][163] = 4'b0111; // x=163, y=34
        pixel_data[34][164] = 4'b0111; // x=164, y=34
        pixel_data[34][165] = 4'b0111; // x=165, y=34
        pixel_data[34][166] = 4'b0111; // x=166, y=34
        pixel_data[34][167] = 4'b0111; // x=167, y=34
        pixel_data[34][168] = 4'b0111; // x=168, y=34
        pixel_data[34][169] = 4'b0111; // x=169, y=34
        pixel_data[34][170] = 4'b0111; // x=170, y=34
        pixel_data[34][171] = 4'b0111; // x=171, y=34
        pixel_data[34][172] = 4'b0111; // x=172, y=34
        pixel_data[34][173] = 4'b0111; // x=173, y=34
        pixel_data[34][174] = 4'b0111; // x=174, y=34
        pixel_data[34][175] = 4'b0111; // x=175, y=34
        pixel_data[34][176] = 4'b0111; // x=176, y=34
        pixel_data[34][177] = 4'b0111; // x=177, y=34
        pixel_data[34][178] = 4'b0111; // x=178, y=34
        pixel_data[34][179] = 4'b0111; // x=179, y=34
        pixel_data[35][0] = 4'b0111; // x=0, y=35
        pixel_data[35][1] = 4'b0111; // x=1, y=35
        pixel_data[35][2] = 4'b0111; // x=2, y=35
        pixel_data[35][3] = 4'b0111; // x=3, y=35
        pixel_data[35][4] = 4'b0111; // x=4, y=35
        pixel_data[35][5] = 4'b0111; // x=5, y=35
        pixel_data[35][6] = 4'b0000; // x=6, y=35
        pixel_data[35][7] = 4'b0000; // x=7, y=35
        pixel_data[35][8] = 4'b0111; // x=8, y=35
        pixel_data[35][9] = 4'b0000; // x=9, y=35
        pixel_data[35][10] = 4'b1111; // x=10, y=35
        pixel_data[35][11] = 4'b1101; // x=11, y=35
        pixel_data[35][12] = 4'b1101; // x=12, y=35
        pixel_data[35][13] = 4'b1100; // x=13, y=35
        pixel_data[35][14] = 4'b0110; // x=14, y=35
        pixel_data[35][15] = 4'b0111; // x=15, y=35
        pixel_data[35][16] = 4'b0000; // x=16, y=35
        pixel_data[35][17] = 4'b0000; // x=17, y=35
        pixel_data[35][18] = 4'b0000; // x=18, y=35
        pixel_data[35][19] = 4'b0000; // x=19, y=35
        pixel_data[35][20] = 4'b0000; // x=20, y=35
        pixel_data[35][21] = 4'b0111; // x=21, y=35
        pixel_data[35][22] = 4'b0000; // x=22, y=35
        pixel_data[35][23] = 4'b0000; // x=23, y=35
        pixel_data[35][24] = 4'b0000; // x=24, y=35
        pixel_data[35][25] = 4'b0111; // x=25, y=35
        pixel_data[35][26] = 4'b1100; // x=26, y=35
        pixel_data[35][27] = 4'b1101; // x=27, y=35
        pixel_data[35][28] = 4'b0001; // x=28, y=35
        pixel_data[35][29] = 4'b0001; // x=29, y=35
        pixel_data[35][30] = 4'b1101; // x=30, y=35
        pixel_data[35][31] = 4'b1000; // x=31, y=35
        pixel_data[35][32] = 4'b0111; // x=32, y=35
        pixel_data[35][33] = 4'b0000; // x=33, y=35
        pixel_data[35][34] = 4'b0000; // x=34, y=35
        pixel_data[35][35] = 4'b0111; // x=35, y=35
        pixel_data[35][36] = 4'b0101; // x=36, y=35
        pixel_data[35][37] = 4'b1101; // x=37, y=35
        pixel_data[35][38] = 4'b0001; // x=38, y=35
        pixel_data[35][39] = 4'b0001; // x=39, y=35
        pixel_data[35][40] = 4'b1101; // x=40, y=35
        pixel_data[35][41] = 4'b1011; // x=41, y=35
        pixel_data[35][42] = 4'b0110; // x=42, y=35
        pixel_data[35][43] = 4'b0111; // x=43, y=35
        pixel_data[35][44] = 4'b0000; // x=44, y=35
        pixel_data[35][45] = 4'b0000; // x=45, y=35
        pixel_data[35][46] = 4'b0000; // x=46, y=35
        pixel_data[35][47] = 4'b0111; // x=47, y=35
        pixel_data[35][48] = 4'b0000; // x=48, y=35
        pixel_data[35][49] = 4'b0000; // x=49, y=35
        pixel_data[35][50] = 4'b0000; // x=50, y=35
        pixel_data[35][51] = 4'b0111; // x=51, y=35
        pixel_data[35][52] = 4'b0111; // x=52, y=35
        pixel_data[35][53] = 4'b0110; // x=53, y=35
        pixel_data[35][54] = 4'b0000; // x=54, y=35
        pixel_data[35][55] = 4'b0111; // x=55, y=35
        pixel_data[35][56] = 4'b0000; // x=56, y=35
        pixel_data[35][57] = 4'b0000; // x=57, y=35
        pixel_data[35][58] = 4'b0111; // x=58, y=35
        pixel_data[35][59] = 4'b0100; // x=59, y=35
        pixel_data[35][60] = 4'b0001; // x=60, y=35
        pixel_data[35][61] = 4'b0001; // x=61, y=35
        pixel_data[35][62] = 4'b1101; // x=62, y=35
        pixel_data[35][63] = 4'b0001; // x=63, y=35
        pixel_data[35][64] = 4'b1101; // x=64, y=35
        pixel_data[35][65] = 4'b1111; // x=65, y=35
        pixel_data[35][66] = 4'b0111; // x=66, y=35
        pixel_data[35][67] = 4'b0111; // x=67, y=35
        pixel_data[35][68] = 4'b0000; // x=68, y=35
        pixel_data[35][69] = 4'b0000; // x=69, y=35
        pixel_data[35][70] = 4'b0111; // x=70, y=35
        pixel_data[35][71] = 4'b0111; // x=71, y=35
        pixel_data[35][72] = 4'b0111; // x=72, y=35
        pixel_data[35][73] = 4'b0000; // x=73, y=35
        pixel_data[35][74] = 4'b0000; // x=74, y=35
        pixel_data[35][75] = 4'b0111; // x=75, y=35
        pixel_data[35][76] = 4'b1010; // x=76, y=35
        pixel_data[35][77] = 4'b1101; // x=77, y=35
        pixel_data[35][78] = 4'b0001; // x=78, y=35
        pixel_data[35][79] = 4'b1101; // x=79, y=35
        pixel_data[35][80] = 4'b0001; // x=80, y=35
        pixel_data[35][81] = 4'b1101; // x=81, y=35
        pixel_data[35][82] = 4'b1010; // x=82, y=35
        pixel_data[35][83] = 4'b0111; // x=83, y=35
        pixel_data[35][84] = 4'b0000; // x=84, y=35
        pixel_data[35][85] = 4'b0000; // x=85, y=35
        pixel_data[35][86] = 4'b0111; // x=86, y=35
        pixel_data[35][87] = 4'b0110; // x=87, y=35
        pixel_data[35][88] = 4'b1011; // x=88, y=35
        pixel_data[35][89] = 4'b1101; // x=89, y=35
        pixel_data[35][90] = 4'b0001; // x=90, y=35
        pixel_data[35][91] = 4'b0001; // x=91, y=35
        pixel_data[35][92] = 4'b1101; // x=92, y=35
        pixel_data[35][93] = 4'b1001; // x=93, y=35
        pixel_data[35][94] = 4'b0111; // x=94, y=35
        pixel_data[35][95] = 4'b0000; // x=95, y=35
        pixel_data[35][96] = 4'b0111; // x=96, y=35
        pixel_data[35][97] = 4'b0111; // x=97, y=35
        pixel_data[35][98] = 4'b0111; // x=98, y=35
        pixel_data[35][99] = 4'b0111; // x=99, y=35
        pixel_data[35][100] = 4'b0111; // x=100, y=35
        pixel_data[35][101] = 4'b0111; // x=101, y=35
        pixel_data[35][102] = 4'b0111; // x=102, y=35
        pixel_data[35][103] = 4'b0111; // x=103, y=35
        pixel_data[35][104] = 4'b1000; // x=104, y=35
        pixel_data[35][105] = 4'b1101; // x=105, y=35
        pixel_data[35][106] = 4'b0001; // x=106, y=35
        pixel_data[35][107] = 4'b1101; // x=107, y=35
        pixel_data[35][108] = 4'b1101; // x=108, y=35
        pixel_data[35][109] = 4'b1011; // x=109, y=35
        pixel_data[35][110] = 4'b0110; // x=110, y=35
        pixel_data[35][111] = 4'b0111; // x=111, y=35
        pixel_data[35][112] = 4'b0000; // x=112, y=35
        pixel_data[35][113] = 4'b0000; // x=113, y=35
        pixel_data[35][114] = 4'b0000; // x=114, y=35
        pixel_data[35][115] = 4'b0000; // x=115, y=35
        pixel_data[35][116] = 4'b0000; // x=116, y=35
        pixel_data[35][117] = 4'b0000; // x=117, y=35
        pixel_data[35][118] = 4'b0000; // x=118, y=35
        pixel_data[35][119] = 4'b0000; // x=119, y=35
        pixel_data[35][120] = 4'b0000; // x=120, y=35
        pixel_data[35][121] = 4'b0111; // x=121, y=35
        pixel_data[35][122] = 4'b0111; // x=122, y=35
        pixel_data[35][123] = 4'b0000; // x=123, y=35
        pixel_data[35][124] = 4'b0000; // x=124, y=35
        pixel_data[35][125] = 4'b0000; // x=125, y=35
        pixel_data[35][126] = 4'b0111; // x=126, y=35
        pixel_data[35][127] = 4'b0111; // x=127, y=35
        pixel_data[35][128] = 4'b0111; // x=128, y=35
        pixel_data[35][129] = 4'b0111; // x=129, y=35
        pixel_data[35][130] = 4'b0111; // x=130, y=35
        pixel_data[35][131] = 4'b0111; // x=131, y=35
        pixel_data[35][132] = 4'b0111; // x=132, y=35
        pixel_data[35][133] = 4'b0111; // x=133, y=35
        pixel_data[35][134] = 4'b0111; // x=134, y=35
        pixel_data[35][135] = 4'b0111; // x=135, y=35
        pixel_data[35][136] = 4'b0111; // x=136, y=35
        pixel_data[35][137] = 4'b0111; // x=137, y=35
        pixel_data[35][138] = 4'b0111; // x=138, y=35
        pixel_data[35][139] = 4'b0111; // x=139, y=35
        pixel_data[35][140] = 4'b0111; // x=140, y=35
        pixel_data[35][141] = 4'b0111; // x=141, y=35
        pixel_data[35][142] = 4'b0000; // x=142, y=35
        pixel_data[35][143] = 4'b0111; // x=143, y=35
        pixel_data[35][144] = 4'b0111; // x=144, y=35
        pixel_data[35][145] = 4'b0111; // x=145, y=35
        pixel_data[35][146] = 4'b0111; // x=146, y=35
        pixel_data[35][147] = 4'b0111; // x=147, y=35
        pixel_data[35][148] = 4'b0111; // x=148, y=35
        pixel_data[35][149] = 4'b0111; // x=149, y=35
        pixel_data[35][150] = 4'b0111; // x=150, y=35
        pixel_data[35][151] = 4'b0111; // x=151, y=35
        pixel_data[35][152] = 4'b0111; // x=152, y=35
        pixel_data[35][153] = 4'b0111; // x=153, y=35
        pixel_data[35][154] = 4'b0111; // x=154, y=35
        pixel_data[35][155] = 4'b0111; // x=155, y=35
        pixel_data[35][156] = 4'b0111; // x=156, y=35
        pixel_data[35][157] = 4'b0111; // x=157, y=35
        pixel_data[35][158] = 4'b0111; // x=158, y=35
        pixel_data[35][159] = 4'b0111; // x=159, y=35
        pixel_data[35][160] = 4'b0111; // x=160, y=35
        pixel_data[35][161] = 4'b0111; // x=161, y=35
        pixel_data[35][162] = 4'b0111; // x=162, y=35
        pixel_data[35][163] = 4'b0111; // x=163, y=35
        pixel_data[35][164] = 4'b0111; // x=164, y=35
        pixel_data[35][165] = 4'b0111; // x=165, y=35
        pixel_data[35][166] = 4'b0111; // x=166, y=35
        pixel_data[35][167] = 4'b0111; // x=167, y=35
        pixel_data[35][168] = 4'b0111; // x=168, y=35
        pixel_data[35][169] = 4'b0111; // x=169, y=35
        pixel_data[35][170] = 4'b0111; // x=170, y=35
        pixel_data[35][171] = 4'b0111; // x=171, y=35
        pixel_data[35][172] = 4'b0111; // x=172, y=35
        pixel_data[35][173] = 4'b0111; // x=173, y=35
        pixel_data[35][174] = 4'b0111; // x=174, y=35
        pixel_data[35][175] = 4'b0111; // x=175, y=35
        pixel_data[35][176] = 4'b0111; // x=176, y=35
        pixel_data[35][177] = 4'b0111; // x=177, y=35
        pixel_data[35][178] = 4'b0111; // x=178, y=35
        pixel_data[35][179] = 4'b0111; // x=179, y=35
        pixel_data[36][0] = 4'b0111; // x=0, y=36
        pixel_data[36][1] = 4'b0111; // x=1, y=36
        pixel_data[36][2] = 4'b0111; // x=2, y=36
        pixel_data[36][3] = 4'b0111; // x=3, y=36
        pixel_data[36][4] = 4'b0111; // x=4, y=36
        pixel_data[36][5] = 4'b0000; // x=5, y=36
        pixel_data[36][6] = 4'b0000; // x=6, y=36
        pixel_data[36][7] = 4'b0000; // x=7, y=36
        pixel_data[36][8] = 4'b0110; // x=8, y=36
        pixel_data[36][9] = 4'b1100; // x=9, y=36
        pixel_data[36][10] = 4'b1101; // x=10, y=36
        pixel_data[36][11] = 4'b0001; // x=11, y=36
        pixel_data[36][12] = 4'b0001; // x=12, y=36
        pixel_data[36][13] = 4'b1101; // x=13, y=36
        pixel_data[36][14] = 4'b1011; // x=14, y=36
        pixel_data[36][15] = 4'b1010; // x=15, y=36
        pixel_data[36][16] = 4'b0000; // x=16, y=36
        pixel_data[36][17] = 4'b0111; // x=17, y=36
        pixel_data[36][18] = 4'b0111; // x=18, y=36
        pixel_data[36][19] = 4'b0111; // x=19, y=36
        pixel_data[36][20] = 4'b0111; // x=20, y=36
        pixel_data[36][21] = 4'b0111; // x=21, y=36
        pixel_data[36][22] = 4'b0111; // x=22, y=36
        pixel_data[36][23] = 4'b0111; // x=23, y=36
        pixel_data[36][24] = 4'b0111; // x=24, y=36
        pixel_data[36][25] = 4'b1010; // x=25, y=36
        pixel_data[36][26] = 4'b1101; // x=26, y=36
        pixel_data[36][27] = 4'b0001; // x=27, y=36
        pixel_data[36][28] = 4'b0001; // x=28, y=36
        pixel_data[36][29] = 4'b0001; // x=29, y=36
        pixel_data[36][30] = 4'b1101; // x=30, y=36
        pixel_data[36][31] = 4'b0010; // x=31, y=36
        pixel_data[36][32] = 4'b0111; // x=32, y=36
        pixel_data[36][33] = 4'b0000; // x=33, y=36
        pixel_data[36][34] = 4'b0111; // x=34, y=36
        pixel_data[36][35] = 4'b0111; // x=35, y=36
        pixel_data[36][36] = 4'b0110; // x=36, y=36
        pixel_data[36][37] = 4'b1011; // x=37, y=36
        pixel_data[36][38] = 4'b1101; // x=38, y=36
        pixel_data[36][39] = 4'b0001; // x=39, y=36
        pixel_data[36][40] = 4'b0001; // x=40, y=36
        pixel_data[36][41] = 4'b1101; // x=41, y=36
        pixel_data[36][42] = 4'b0011; // x=42, y=36
        pixel_data[36][43] = 4'b0100; // x=43, y=36
        pixel_data[36][44] = 4'b0111; // x=44, y=36
        pixel_data[36][45] = 4'b0111; // x=45, y=36
        pixel_data[36][46] = 4'b0111; // x=46, y=36
        pixel_data[36][47] = 4'b0111; // x=47, y=36
        pixel_data[36][48] = 4'b0111; // x=48, y=36
        pixel_data[36][49] = 4'b0111; // x=49, y=36
        pixel_data[36][50] = 4'b0111; // x=50, y=36
        pixel_data[36][51] = 4'b0000; // x=51, y=36
        pixel_data[36][52] = 4'b0010; // x=52, y=36
        pixel_data[36][53] = 4'b0001; // x=53, y=36
        pixel_data[36][54] = 4'b1111; // x=54, y=36
        pixel_data[36][55] = 4'b0000; // x=55, y=36
        pixel_data[36][56] = 4'b0111; // x=56, y=36
        pixel_data[36][57] = 4'b0000; // x=57, y=36
        pixel_data[36][58] = 4'b0000; // x=58, y=36
        pixel_data[36][59] = 4'b0111; // x=59, y=36
        pixel_data[36][60] = 4'b1111; // x=60, y=36
        pixel_data[36][61] = 4'b1101; // x=61, y=36
        pixel_data[36][62] = 4'b0001; // x=62, y=36
        pixel_data[36][63] = 4'b0001; // x=63, y=36
        pixel_data[36][64] = 4'b0001; // x=64, y=36
        pixel_data[36][65] = 4'b1101; // x=65, y=36
        pixel_data[36][66] = 4'b0101; // x=66, y=36
        pixel_data[36][67] = 4'b0000; // x=67, y=36
        pixel_data[36][68] = 4'b0111; // x=68, y=36
        pixel_data[36][69] = 4'b0111; // x=69, y=36
        pixel_data[36][70] = 4'b0111; // x=70, y=36
        pixel_data[36][71] = 4'b0111; // x=71, y=36
        pixel_data[36][72] = 4'b0111; // x=72, y=36
        pixel_data[36][73] = 4'b0111; // x=73, y=36
        pixel_data[36][74] = 4'b0111; // x=74, y=36
        pixel_data[36][75] = 4'b1010; // x=75, y=36
        pixel_data[36][76] = 4'b0001; // x=76, y=36
        pixel_data[36][77] = 4'b1101; // x=77, y=36
        pixel_data[36][78] = 4'b1101; // x=78, y=36
        pixel_data[36][79] = 4'b0001; // x=79, y=36
        pixel_data[36][80] = 4'b1101; // x=80, y=36
        pixel_data[36][81] = 4'b0011; // x=81, y=36
        pixel_data[36][82] = 4'b0000; // x=82, y=36
        pixel_data[36][83] = 4'b0111; // x=83, y=36
        pixel_data[36][84] = 4'b0000; // x=84, y=36
        pixel_data[36][85] = 4'b0111; // x=85, y=36
        pixel_data[36][86] = 4'b0111; // x=86, y=36
        pixel_data[36][87] = 4'b0110; // x=87, y=36
        pixel_data[36][88] = 4'b1011; // x=88, y=36
        pixel_data[36][89] = 4'b1101; // x=89, y=36
        pixel_data[36][90] = 4'b0001; // x=90, y=36
        pixel_data[36][91] = 4'b0001; // x=91, y=36
        pixel_data[36][92] = 4'b1101; // x=92, y=36
        pixel_data[36][93] = 4'b1001; // x=93, y=36
        pixel_data[36][94] = 4'b0111; // x=94, y=36
        pixel_data[36][95] = 4'b0000; // x=95, y=36
        pixel_data[36][96] = 4'b0111; // x=96, y=36
        pixel_data[36][97] = 4'b0111; // x=97, y=36
        pixel_data[36][98] = 4'b0111; // x=98, y=36
        pixel_data[36][99] = 4'b0111; // x=99, y=36
        pixel_data[36][100] = 4'b0111; // x=100, y=36
        pixel_data[36][101] = 4'b0111; // x=101, y=36
        pixel_data[36][102] = 4'b0111; // x=102, y=36
        pixel_data[36][103] = 4'b0111; // x=103, y=36
        pixel_data[36][104] = 4'b0100; // x=104, y=36
        pixel_data[36][105] = 4'b0001; // x=105, y=36
        pixel_data[36][106] = 4'b0001; // x=106, y=36
        pixel_data[36][107] = 4'b0001; // x=107, y=36
        pixel_data[36][108] = 4'b0001; // x=108, y=36
        pixel_data[36][109] = 4'b1101; // x=109, y=36
        pixel_data[36][110] = 4'b0011; // x=110, y=36
        pixel_data[36][111] = 4'b0100; // x=111, y=36
        pixel_data[36][112] = 4'b0111; // x=112, y=36
        pixel_data[36][113] = 4'b0111; // x=113, y=36
        pixel_data[36][114] = 4'b0111; // x=114, y=36
        pixel_data[36][115] = 4'b0111; // x=115, y=36
        pixel_data[36][116] = 4'b0111; // x=116, y=36
        pixel_data[36][117] = 4'b0111; // x=117, y=36
        pixel_data[36][118] = 4'b0111; // x=118, y=36
        pixel_data[36][119] = 4'b0111; // x=119, y=36
        pixel_data[36][120] = 4'b0111; // x=120, y=36
        pixel_data[36][121] = 4'b1001; // x=121, y=36
        pixel_data[36][122] = 4'b0101; // x=122, y=36
        pixel_data[36][123] = 4'b0000; // x=123, y=36
        pixel_data[36][124] = 4'b0000; // x=124, y=36
        pixel_data[36][125] = 4'b0000; // x=125, y=36
        pixel_data[36][126] = 4'b0111; // x=126, y=36
        pixel_data[36][127] = 4'b0111; // x=127, y=36
        pixel_data[36][128] = 4'b0111; // x=128, y=36
        pixel_data[36][129] = 4'b0111; // x=129, y=36
        pixel_data[36][130] = 4'b0111; // x=130, y=36
        pixel_data[36][131] = 4'b0111; // x=131, y=36
        pixel_data[36][132] = 4'b0111; // x=132, y=36
        pixel_data[36][133] = 4'b0111; // x=133, y=36
        pixel_data[36][134] = 4'b0111; // x=134, y=36
        pixel_data[36][135] = 4'b0111; // x=135, y=36
        pixel_data[36][136] = 4'b0111; // x=136, y=36
        pixel_data[36][137] = 4'b0111; // x=137, y=36
        pixel_data[36][138] = 4'b0111; // x=138, y=36
        pixel_data[36][139] = 4'b0111; // x=139, y=36
        pixel_data[36][140] = 4'b0111; // x=140, y=36
        pixel_data[36][141] = 4'b0000; // x=141, y=36
        pixel_data[36][142] = 4'b0111; // x=142, y=36
        pixel_data[36][143] = 4'b1110; // x=143, y=36
        pixel_data[36][144] = 4'b0010; // x=144, y=36
        pixel_data[36][145] = 4'b1111; // x=145, y=36
        pixel_data[36][146] = 4'b0101; // x=146, y=36
        pixel_data[36][147] = 4'b0100; // x=147, y=36
        pixel_data[36][148] = 4'b0111; // x=148, y=36
        pixel_data[36][149] = 4'b0000; // x=149, y=36
        pixel_data[36][150] = 4'b0111; // x=150, y=36
        pixel_data[36][151] = 4'b0000; // x=151, y=36
        pixel_data[36][152] = 4'b0111; // x=152, y=36
        pixel_data[36][153] = 4'b0111; // x=153, y=36
        pixel_data[36][154] = 4'b0111; // x=154, y=36
        pixel_data[36][155] = 4'b0111; // x=155, y=36
        pixel_data[36][156] = 4'b0111; // x=156, y=36
        pixel_data[36][157] = 4'b0111; // x=157, y=36
        pixel_data[36][158] = 4'b0111; // x=158, y=36
        pixel_data[36][159] = 4'b0111; // x=159, y=36
        pixel_data[36][160] = 4'b0111; // x=160, y=36
        pixel_data[36][161] = 4'b0111; // x=161, y=36
        pixel_data[36][162] = 4'b0111; // x=162, y=36
        pixel_data[36][163] = 4'b0111; // x=163, y=36
        pixel_data[36][164] = 4'b0111; // x=164, y=36
        pixel_data[36][165] = 4'b0111; // x=165, y=36
        pixel_data[36][166] = 4'b0111; // x=166, y=36
        pixel_data[36][167] = 4'b0111; // x=167, y=36
        pixel_data[36][168] = 4'b0111; // x=168, y=36
        pixel_data[36][169] = 4'b0111; // x=169, y=36
        pixel_data[36][170] = 4'b0111; // x=170, y=36
        pixel_data[36][171] = 4'b0111; // x=171, y=36
        pixel_data[36][172] = 4'b0111; // x=172, y=36
        pixel_data[36][173] = 4'b0111; // x=173, y=36
        pixel_data[36][174] = 4'b0111; // x=174, y=36
        pixel_data[36][175] = 4'b0111; // x=175, y=36
        pixel_data[36][176] = 4'b0111; // x=176, y=36
        pixel_data[36][177] = 4'b0111; // x=177, y=36
        pixel_data[36][178] = 4'b0111; // x=178, y=36
        pixel_data[36][179] = 4'b0111; // x=179, y=36
        pixel_data[37][0] = 4'b0111; // x=0, y=37
        pixel_data[37][1] = 4'b0111; // x=1, y=37
        pixel_data[37][2] = 4'b0111; // x=2, y=37
        pixel_data[37][3] = 4'b0111; // x=3, y=37
        pixel_data[37][4] = 4'b0111; // x=4, y=37
        pixel_data[37][5] = 4'b0000; // x=5, y=37
        pixel_data[37][6] = 4'b0000; // x=6, y=37
        pixel_data[37][7] = 4'b0111; // x=7, y=37
        pixel_data[37][8] = 4'b0100; // x=8, y=37
        pixel_data[37][9] = 4'b1011; // x=9, y=37
        pixel_data[37][10] = 4'b1101; // x=10, y=37
        pixel_data[37][11] = 4'b0001; // x=11, y=37
        pixel_data[37][12] = 4'b1101; // x=12, y=37
        pixel_data[37][13] = 4'b0001; // x=13, y=37
        pixel_data[37][14] = 4'b1101; // x=14, y=37
        pixel_data[37][15] = 4'b1101; // x=15, y=37
        pixel_data[37][16] = 4'b0011; // x=16, y=37
        pixel_data[37][17] = 4'b0101; // x=17, y=37
        pixel_data[37][18] = 4'b1001; // x=18, y=37
        pixel_data[37][19] = 4'b0100; // x=19, y=37
        pixel_data[37][20] = 4'b0110; // x=20, y=37
        pixel_data[37][21] = 4'b1110; // x=21, y=37
        pixel_data[37][22] = 4'b0100; // x=22, y=37
        pixel_data[37][23] = 4'b1010; // x=23, y=37
        pixel_data[37][24] = 4'b1100; // x=24, y=37
        pixel_data[37][25] = 4'b1101; // x=25, y=37
        pixel_data[37][26] = 4'b0001; // x=26, y=37
        pixel_data[37][27] = 4'b1101; // x=27, y=37
        pixel_data[37][28] = 4'b0001; // x=28, y=37
        pixel_data[37][29] = 4'b1101; // x=29, y=37
        pixel_data[37][30] = 4'b1011; // x=30, y=37
        pixel_data[37][31] = 4'b1110; // x=31, y=37
        pixel_data[37][32] = 4'b0111; // x=32, y=37
        pixel_data[37][33] = 4'b0111; // x=33, y=37
        pixel_data[37][34] = 4'b0111; // x=34, y=37
        pixel_data[37][35] = 4'b0000; // x=35, y=37
        pixel_data[37][36] = 4'b0111; // x=36, y=37
        pixel_data[37][37] = 4'b0010; // x=37, y=37
        pixel_data[37][38] = 4'b1101; // x=38, y=37
        pixel_data[37][39] = 4'b0001; // x=39, y=37
        pixel_data[37][40] = 4'b0001; // x=40, y=37
        pixel_data[37][41] = 4'b0001; // x=41, y=37
        pixel_data[37][42] = 4'b1101; // x=42, y=37
        pixel_data[37][43] = 4'b1101; // x=43, y=37
        pixel_data[37][44] = 4'b1111; // x=44, y=37
        pixel_data[37][45] = 4'b0100; // x=45, y=37
        pixel_data[37][46] = 4'b1110; // x=46, y=37
        pixel_data[37][47] = 4'b1110; // x=47, y=37
        pixel_data[37][48] = 4'b1110; // x=48, y=37
        pixel_data[37][49] = 4'b0110; // x=49, y=37
        pixel_data[37][50] = 4'b1010; // x=50, y=37
        pixel_data[37][51] = 4'b0011; // x=51, y=37
        pixel_data[37][52] = 4'b1101; // x=52, y=37
        pixel_data[37][53] = 4'b0001; // x=53, y=37
        pixel_data[37][54] = 4'b1101; // x=54, y=37
        pixel_data[37][55] = 4'b1111; // x=55, y=37
        pixel_data[37][56] = 4'b1110; // x=56, y=37
        pixel_data[37][57] = 4'b0000; // x=57, y=37
        pixel_data[37][58] = 4'b0000; // x=58, y=37
        pixel_data[37][59] = 4'b0111; // x=59, y=37
        pixel_data[37][60] = 4'b0110; // x=60, y=37
        pixel_data[37][61] = 4'b1011; // x=61, y=37
        pixel_data[37][62] = 4'b1101; // x=62, y=37
        pixel_data[37][63] = 4'b0001; // x=63, y=37
        pixel_data[37][64] = 4'b0001; // x=64, y=37
        pixel_data[37][65] = 4'b0001; // x=65, y=37
        pixel_data[37][66] = 4'b1101; // x=66, y=37
        pixel_data[37][67] = 4'b1100; // x=67, y=37
        pixel_data[37][68] = 4'b1010; // x=68, y=37
        pixel_data[37][69] = 4'b0110; // x=69, y=37
        pixel_data[37][70] = 4'b1110; // x=70, y=37
        pixel_data[37][71] = 4'b1110; // x=71, y=37
        pixel_data[37][72] = 4'b1110; // x=72, y=37
        pixel_data[37][73] = 4'b1001; // x=73, y=37
        pixel_data[37][74] = 4'b1000; // x=74, y=37
        pixel_data[37][75] = 4'b1101; // x=75, y=37
        pixel_data[37][76] = 4'b0001; // x=76, y=37
        pixel_data[37][77] = 4'b1101; // x=77, y=37
        pixel_data[37][78] = 4'b0001; // x=78, y=37
        pixel_data[37][79] = 4'b0001; // x=79, y=37
        pixel_data[37][80] = 4'b0001; // x=80, y=37
        pixel_data[37][81] = 4'b0100; // x=81, y=37
        pixel_data[37][82] = 4'b0111; // x=82, y=37
        pixel_data[37][83] = 4'b0000; // x=83, y=37
        pixel_data[37][84] = 4'b0111; // x=84, y=37
        pixel_data[37][85] = 4'b0000; // x=85, y=37
        pixel_data[37][86] = 4'b0111; // x=86, y=37
        pixel_data[37][87] = 4'b0110; // x=87, y=37
        pixel_data[37][88] = 4'b1011; // x=88, y=37
        pixel_data[37][89] = 4'b1101; // x=89, y=37
        pixel_data[37][90] = 4'b0001; // x=90, y=37
        pixel_data[37][91] = 4'b0001; // x=91, y=37
        pixel_data[37][92] = 4'b1101; // x=92, y=37
        pixel_data[37][93] = 4'b1001; // x=93, y=37
        pixel_data[37][94] = 4'b0111; // x=94, y=37
        pixel_data[37][95] = 4'b0000; // x=95, y=37
        pixel_data[37][96] = 4'b0111; // x=96, y=37
        pixel_data[37][97] = 4'b0111; // x=97, y=37
        pixel_data[37][98] = 4'b0111; // x=98, y=37
        pixel_data[37][99] = 4'b0111; // x=99, y=37
        pixel_data[37][100] = 4'b0111; // x=100, y=37
        pixel_data[37][101] = 4'b0111; // x=101, y=37
        pixel_data[37][102] = 4'b0111; // x=102, y=37
        pixel_data[37][103] = 4'b0000; // x=103, y=37
        pixel_data[37][104] = 4'b0111; // x=104, y=37
        pixel_data[37][105] = 4'b0101; // x=105, y=37
        pixel_data[37][106] = 4'b1101; // x=106, y=37
        pixel_data[37][107] = 4'b0001; // x=107, y=37
        pixel_data[37][108] = 4'b0001; // x=108, y=37
        pixel_data[37][109] = 4'b0001; // x=109, y=37
        pixel_data[37][110] = 4'b1101; // x=110, y=37
        pixel_data[37][111] = 4'b1101; // x=111, y=37
        pixel_data[37][112] = 4'b1111; // x=112, y=37
        pixel_data[37][113] = 4'b1010; // x=113, y=37
        pixel_data[37][114] = 4'b0110; // x=114, y=37
        pixel_data[37][115] = 4'b1110; // x=115, y=37
        pixel_data[37][116] = 4'b1110; // x=116, y=37
        pixel_data[37][117] = 4'b1110; // x=117, y=37
        pixel_data[37][118] = 4'b0110; // x=118, y=37
        pixel_data[37][119] = 4'b1010; // x=119, y=37
        pixel_data[37][120] = 4'b1100; // x=120, y=37
        pixel_data[37][121] = 4'b1101; // x=121, y=37
        pixel_data[37][122] = 4'b1101; // x=122, y=37
        pixel_data[37][123] = 4'b1111; // x=123, y=37
        pixel_data[37][124] = 4'b0111; // x=124, y=37
        pixel_data[37][125] = 4'b0000; // x=125, y=37
        pixel_data[37][126] = 4'b0111; // x=126, y=37
        pixel_data[37][127] = 4'b0111; // x=127, y=37
        pixel_data[37][128] = 4'b0111; // x=128, y=37
        pixel_data[37][129] = 4'b0111; // x=129, y=37
        pixel_data[37][130] = 4'b0111; // x=130, y=37
        pixel_data[37][131] = 4'b0111; // x=131, y=37
        pixel_data[37][132] = 4'b0111; // x=132, y=37
        pixel_data[37][133] = 4'b0111; // x=133, y=37
        pixel_data[37][134] = 4'b0111; // x=134, y=37
        pixel_data[37][135] = 4'b0111; // x=135, y=37
        pixel_data[37][136] = 4'b0111; // x=136, y=37
        pixel_data[37][137] = 4'b0111; // x=137, y=37
        pixel_data[37][138] = 4'b0111; // x=138, y=37
        pixel_data[37][139] = 4'b0111; // x=139, y=37
        pixel_data[37][140] = 4'b0000; // x=140, y=37
        pixel_data[37][141] = 4'b0111; // x=141, y=37
        pixel_data[37][142] = 4'b1110; // x=142, y=37
        pixel_data[37][143] = 4'b0011; // x=143, y=37
        pixel_data[37][144] = 4'b1101; // x=144, y=37
        pixel_data[37][145] = 4'b1101; // x=145, y=37
        pixel_data[37][146] = 4'b1101; // x=146, y=37
        pixel_data[37][147] = 4'b1101; // x=147, y=37
        pixel_data[37][148] = 4'b1010; // x=148, y=37
        pixel_data[37][149] = 4'b0111; // x=149, y=37
        pixel_data[37][150] = 4'b0000; // x=150, y=37
        pixel_data[37][151] = 4'b0000; // x=151, y=37
        pixel_data[37][152] = 4'b0111; // x=152, y=37
        pixel_data[37][153] = 4'b0111; // x=153, y=37
        pixel_data[37][154] = 4'b0111; // x=154, y=37
        pixel_data[37][155] = 4'b0111; // x=155, y=37
        pixel_data[37][156] = 4'b0111; // x=156, y=37
        pixel_data[37][157] = 4'b0111; // x=157, y=37
        pixel_data[37][158] = 4'b0111; // x=158, y=37
        pixel_data[37][159] = 4'b0111; // x=159, y=37
        pixel_data[37][160] = 4'b0111; // x=160, y=37
        pixel_data[37][161] = 4'b0111; // x=161, y=37
        pixel_data[37][162] = 4'b0111; // x=162, y=37
        pixel_data[37][163] = 4'b0111; // x=163, y=37
        pixel_data[37][164] = 4'b0111; // x=164, y=37
        pixel_data[37][165] = 4'b0111; // x=165, y=37
        pixel_data[37][166] = 4'b0111; // x=166, y=37
        pixel_data[37][167] = 4'b0111; // x=167, y=37
        pixel_data[37][168] = 4'b0111; // x=168, y=37
        pixel_data[37][169] = 4'b0111; // x=169, y=37
        pixel_data[37][170] = 4'b0111; // x=170, y=37
        pixel_data[37][171] = 4'b0111; // x=171, y=37
        pixel_data[37][172] = 4'b0111; // x=172, y=37
        pixel_data[37][173] = 4'b0111; // x=173, y=37
        pixel_data[37][174] = 4'b0111; // x=174, y=37
        pixel_data[37][175] = 4'b0111; // x=175, y=37
        pixel_data[37][176] = 4'b0111; // x=176, y=37
        pixel_data[37][177] = 4'b0111; // x=177, y=37
        pixel_data[37][178] = 4'b0111; // x=178, y=37
        pixel_data[37][179] = 4'b0111; // x=179, y=37
        pixel_data[38][0] = 4'b0111; // x=0, y=38
        pixel_data[38][1] = 4'b0111; // x=1, y=38
        pixel_data[38][2] = 4'b0111; // x=2, y=38
        pixel_data[38][3] = 4'b0111; // x=3, y=38
        pixel_data[38][4] = 4'b0111; // x=4, y=38
        pixel_data[38][5] = 4'b0111; // x=5, y=38
        pixel_data[38][6] = 4'b0111; // x=6, y=38
        pixel_data[38][7] = 4'b0000; // x=7, y=38
        pixel_data[38][8] = 4'b0111; // x=8, y=38
        pixel_data[38][9] = 4'b0110; // x=9, y=38
        pixel_data[38][10] = 4'b0011; // x=10, y=38
        pixel_data[38][11] = 4'b1101; // x=11, y=38
        pixel_data[38][12] = 4'b0001; // x=12, y=38
        pixel_data[38][13] = 4'b0001; // x=13, y=38
        pixel_data[38][14] = 4'b0001; // x=14, y=38
        pixel_data[38][15] = 4'b0001; // x=15, y=38
        pixel_data[38][16] = 4'b1101; // x=16, y=38
        pixel_data[38][17] = 4'b1101; // x=17, y=38
        pixel_data[38][18] = 4'b1101; // x=18, y=38
        pixel_data[38][19] = 4'b1101; // x=19, y=38
        pixel_data[38][20] = 4'b0001; // x=20, y=38
        pixel_data[38][21] = 4'b0001; // x=21, y=38
        pixel_data[38][22] = 4'b0001; // x=22, y=38
        pixel_data[38][23] = 4'b1101; // x=23, y=38
        pixel_data[38][24] = 4'b1101; // x=24, y=38
        pixel_data[38][25] = 4'b0001; // x=25, y=38
        pixel_data[38][26] = 4'b0001; // x=26, y=38
        pixel_data[38][27] = 4'b0001; // x=27, y=38
        pixel_data[38][28] = 4'b1101; // x=28, y=38
        pixel_data[38][29] = 4'b0001; // x=29, y=38
        pixel_data[38][30] = 4'b1001; // x=30, y=38
        pixel_data[38][31] = 4'b0111; // x=31, y=38
        pixel_data[38][32] = 4'b0000; // x=32, y=38
        pixel_data[38][33] = 4'b0000; // x=33, y=38
        pixel_data[38][34] = 4'b0111; // x=34, y=38
        pixel_data[38][35] = 4'b0000; // x=35, y=38
        pixel_data[38][36] = 4'b0000; // x=36, y=38
        pixel_data[38][37] = 4'b0111; // x=37, y=38
        pixel_data[38][38] = 4'b0010; // x=38, y=38
        pixel_data[38][39] = 4'b1101; // x=39, y=38
        pixel_data[38][40] = 4'b1101; // x=40, y=38
        pixel_data[38][41] = 4'b0001; // x=41, y=38
        pixel_data[38][42] = 4'b0001; // x=42, y=38
        pixel_data[38][43] = 4'b0001; // x=43, y=38
        pixel_data[38][44] = 4'b1101; // x=44, y=38
        pixel_data[38][45] = 4'b1101; // x=45, y=38
        pixel_data[38][46] = 4'b1011; // x=46, y=38
        pixel_data[38][47] = 4'b0011; // x=47, y=38
        pixel_data[38][48] = 4'b1011; // x=48, y=38
        pixel_data[38][49] = 4'b0001; // x=49, y=38
        pixel_data[38][50] = 4'b1101; // x=50, y=38
        pixel_data[38][51] = 4'b1101; // x=51, y=38
        pixel_data[38][52] = 4'b0001; // x=52, y=38
        pixel_data[38][53] = 4'b0001; // x=53, y=38
        pixel_data[38][54] = 4'b1101; // x=54, y=38
        pixel_data[38][55] = 4'b1101; // x=55, y=38
        pixel_data[38][56] = 4'b1001; // x=56, y=38
        pixel_data[38][57] = 4'b0111; // x=57, y=38
        pixel_data[38][58] = 4'b0000; // x=58, y=38
        pixel_data[38][59] = 4'b0000; // x=59, y=38
        pixel_data[38][60] = 4'b0111; // x=60, y=38
        pixel_data[38][61] = 4'b0100; // x=61, y=38
        pixel_data[38][62] = 4'b1011; // x=62, y=38
        pixel_data[38][63] = 4'b1101; // x=63, y=38
        pixel_data[38][64] = 4'b0001; // x=64, y=38
        pixel_data[38][65] = 4'b0001; // x=65, y=38
        pixel_data[38][66] = 4'b0001; // x=66, y=38
        pixel_data[38][67] = 4'b1101; // x=67, y=38
        pixel_data[38][68] = 4'b1101; // x=68, y=38
        pixel_data[38][69] = 4'b0001; // x=69, y=38
        pixel_data[38][70] = 4'b1011; // x=70, y=38
        pixel_data[38][71] = 4'b1011; // x=71, y=38
        pixel_data[38][72] = 4'b0001; // x=72, y=38
        pixel_data[38][73] = 4'b1101; // x=73, y=38
        pixel_data[38][74] = 4'b1101; // x=74, y=38
        pixel_data[38][75] = 4'b0001; // x=75, y=38
        pixel_data[38][76] = 4'b0001; // x=76, y=38
        pixel_data[38][77] = 4'b0001; // x=77, y=38
        pixel_data[38][78] = 4'b1101; // x=78, y=38
        pixel_data[38][79] = 4'b0001; // x=79, y=38
        pixel_data[38][80] = 4'b1001; // x=80, y=38
        pixel_data[38][81] = 4'b0111; // x=81, y=38
        pixel_data[38][82] = 4'b0000; // x=82, y=38
        pixel_data[38][83] = 4'b0111; // x=83, y=38
        pixel_data[38][84] = 4'b0111; // x=84, y=38
        pixel_data[38][85] = 4'b0000; // x=85, y=38
        pixel_data[38][86] = 4'b0111; // x=86, y=38
        pixel_data[38][87] = 4'b0110; // x=87, y=38
        pixel_data[38][88] = 4'b1011; // x=88, y=38
        pixel_data[38][89] = 4'b1101; // x=89, y=38
        pixel_data[38][90] = 4'b0001; // x=90, y=38
        pixel_data[38][91] = 4'b0001; // x=91, y=38
        pixel_data[38][92] = 4'b1101; // x=92, y=38
        pixel_data[38][93] = 4'b1001; // x=93, y=38
        pixel_data[38][94] = 4'b0111; // x=94, y=38
        pixel_data[38][95] = 4'b0000; // x=95, y=38
        pixel_data[38][96] = 4'b0111; // x=96, y=38
        pixel_data[38][97] = 4'b0111; // x=97, y=38
        pixel_data[38][98] = 4'b0111; // x=98, y=38
        pixel_data[38][99] = 4'b0111; // x=99, y=38
        pixel_data[38][100] = 4'b0111; // x=100, y=38
        pixel_data[38][101] = 4'b0111; // x=101, y=38
        pixel_data[38][102] = 4'b0111; // x=102, y=38
        pixel_data[38][103] = 4'b0111; // x=103, y=38
        pixel_data[38][104] = 4'b0000; // x=104, y=38
        pixel_data[38][105] = 4'b0111; // x=105, y=38
        pixel_data[38][106] = 4'b0101; // x=106, y=38
        pixel_data[38][107] = 4'b1101; // x=107, y=38
        pixel_data[38][108] = 4'b1101; // x=108, y=38
        pixel_data[38][109] = 4'b0001; // x=109, y=38
        pixel_data[38][110] = 4'b0001; // x=110, y=38
        pixel_data[38][111] = 4'b1101; // x=111, y=38
        pixel_data[38][112] = 4'b1101; // x=112, y=38
        pixel_data[38][113] = 4'b1101; // x=113, y=38
        pixel_data[38][114] = 4'b1101; // x=114, y=38
        pixel_data[38][115] = 4'b0001; // x=115, y=38
        pixel_data[38][116] = 4'b1011; // x=116, y=38
        pixel_data[38][117] = 4'b1011; // x=117, y=38
        pixel_data[38][118] = 4'b1101; // x=118, y=38
        pixel_data[38][119] = 4'b1101; // x=119, y=38
        pixel_data[38][120] = 4'b1101; // x=120, y=38
        pixel_data[38][121] = 4'b0001; // x=121, y=38
        pixel_data[38][122] = 4'b1011; // x=122, y=38
        pixel_data[38][123] = 4'b1101; // x=123, y=38
        pixel_data[38][124] = 4'b0101; // x=124, y=38
        pixel_data[38][125] = 4'b0111; // x=125, y=38
        pixel_data[38][126] = 4'b0111; // x=126, y=38
        pixel_data[38][127] = 4'b0111; // x=127, y=38
        pixel_data[38][128] = 4'b0111; // x=128, y=38
        pixel_data[38][129] = 4'b0111; // x=129, y=38
        pixel_data[38][130] = 4'b0111; // x=130, y=38
        pixel_data[38][131] = 4'b0111; // x=131, y=38
        pixel_data[38][132] = 4'b0111; // x=132, y=38
        pixel_data[38][133] = 4'b0111; // x=133, y=38
        pixel_data[38][134] = 4'b0111; // x=134, y=38
        pixel_data[38][135] = 4'b0111; // x=135, y=38
        pixel_data[38][136] = 4'b0111; // x=136, y=38
        pixel_data[38][137] = 4'b0111; // x=137, y=38
        pixel_data[38][138] = 4'b0111; // x=138, y=38
        pixel_data[38][139] = 4'b0111; // x=139, y=38
        pixel_data[38][140] = 4'b0000; // x=140, y=38
        pixel_data[38][141] = 4'b0111; // x=141, y=38
        pixel_data[38][142] = 4'b0010; // x=142, y=38
        pixel_data[38][143] = 4'b1101; // x=143, y=38
        pixel_data[38][144] = 4'b0001; // x=144, y=38
        pixel_data[38][145] = 4'b0001; // x=145, y=38
        pixel_data[38][146] = 4'b0001; // x=146, y=38
        pixel_data[38][147] = 4'b1101; // x=147, y=38
        pixel_data[38][148] = 4'b0011; // x=148, y=38
        pixel_data[38][149] = 4'b0000; // x=149, y=38
        pixel_data[38][150] = 4'b0111; // x=150, y=38
        pixel_data[38][151] = 4'b0000; // x=151, y=38
        pixel_data[38][152] = 4'b0111; // x=152, y=38
        pixel_data[38][153] = 4'b0111; // x=153, y=38
        pixel_data[38][154] = 4'b0111; // x=154, y=38
        pixel_data[38][155] = 4'b0111; // x=155, y=38
        pixel_data[38][156] = 4'b0111; // x=156, y=38
        pixel_data[38][157] = 4'b0111; // x=157, y=38
        pixel_data[38][158] = 4'b0111; // x=158, y=38
        pixel_data[38][159] = 4'b0111; // x=159, y=38
        pixel_data[38][160] = 4'b0111; // x=160, y=38
        pixel_data[38][161] = 4'b0111; // x=161, y=38
        pixel_data[38][162] = 4'b0111; // x=162, y=38
        pixel_data[38][163] = 4'b0111; // x=163, y=38
        pixel_data[38][164] = 4'b0111; // x=164, y=38
        pixel_data[38][165] = 4'b0111; // x=165, y=38
        pixel_data[38][166] = 4'b0111; // x=166, y=38
        pixel_data[38][167] = 4'b0111; // x=167, y=38
        pixel_data[38][168] = 4'b0111; // x=168, y=38
        pixel_data[38][169] = 4'b0111; // x=169, y=38
        pixel_data[38][170] = 4'b0111; // x=170, y=38
        pixel_data[38][171] = 4'b0111; // x=171, y=38
        pixel_data[38][172] = 4'b0111; // x=172, y=38
        pixel_data[38][173] = 4'b0111; // x=173, y=38
        pixel_data[38][174] = 4'b0111; // x=174, y=38
        pixel_data[38][175] = 4'b0111; // x=175, y=38
        pixel_data[38][176] = 4'b0111; // x=176, y=38
        pixel_data[38][177] = 4'b0111; // x=177, y=38
        pixel_data[38][178] = 4'b0111; // x=178, y=38
        pixel_data[38][179] = 4'b0111; // x=179, y=38
        pixel_data[39][0] = 4'b0111; // x=0, y=39
        pixel_data[39][1] = 4'b0111; // x=1, y=39
        pixel_data[39][2] = 4'b0111; // x=2, y=39
        pixel_data[39][3] = 4'b0111; // x=3, y=39
        pixel_data[39][4] = 4'b0111; // x=4, y=39
        pixel_data[39][5] = 4'b0111; // x=5, y=39
        pixel_data[39][6] = 4'b0111; // x=6, y=39
        pixel_data[39][7] = 4'b0111; // x=7, y=39
        pixel_data[39][8] = 4'b0111; // x=8, y=39
        pixel_data[39][9] = 4'b0111; // x=9, y=39
        pixel_data[39][10] = 4'b1110; // x=10, y=39
        pixel_data[39][11] = 4'b0101; // x=11, y=39
        pixel_data[39][12] = 4'b0001; // x=12, y=39
        pixel_data[39][13] = 4'b1101; // x=13, y=39
        pixel_data[39][14] = 4'b1101; // x=14, y=39
        pixel_data[39][15] = 4'b1101; // x=15, y=39
        pixel_data[39][16] = 4'b0001; // x=16, y=39
        pixel_data[39][17] = 4'b0001; // x=17, y=39
        pixel_data[39][18] = 4'b0001; // x=18, y=39
        pixel_data[39][19] = 4'b1101; // x=19, y=39
        pixel_data[39][20] = 4'b1101; // x=20, y=39
        pixel_data[39][21] = 4'b1101; // x=21, y=39
        pixel_data[39][22] = 4'b0001; // x=22, y=39
        pixel_data[39][23] = 4'b0001; // x=23, y=39
        pixel_data[39][24] = 4'b0001; // x=24, y=39
        pixel_data[39][25] = 4'b1101; // x=25, y=39
        pixel_data[39][26] = 4'b1101; // x=26, y=39
        pixel_data[39][27] = 4'b1101; // x=27, y=39
        pixel_data[39][28] = 4'b0011; // x=28, y=39
        pixel_data[39][29] = 4'b0100; // x=29, y=39
        pixel_data[39][30] = 4'b0111; // x=30, y=39
        pixel_data[39][31] = 4'b0000; // x=31, y=39
        pixel_data[39][32] = 4'b0111; // x=32, y=39
        pixel_data[39][33] = 4'b0111; // x=33, y=39
        pixel_data[39][34] = 4'b0111; // x=34, y=39
        pixel_data[39][35] = 4'b0111; // x=35, y=39
        pixel_data[39][36] = 4'b0111; // x=36, y=39
        pixel_data[39][37] = 4'b0000; // x=37, y=39
        pixel_data[39][38] = 4'b0111; // x=38, y=39
        pixel_data[39][39] = 4'b1010; // x=39, y=39
        pixel_data[39][40] = 4'b1011; // x=40, y=39
        pixel_data[39][41] = 4'b1101; // x=41, y=39
        pixel_data[39][42] = 4'b1101; // x=42, y=39
        pixel_data[39][43] = 4'b0001; // x=43, y=39
        pixel_data[39][44] = 4'b0001; // x=44, y=39
        pixel_data[39][45] = 4'b0001; // x=45, y=39
        pixel_data[39][46] = 4'b1101; // x=46, y=39
        pixel_data[39][47] = 4'b1101; // x=47, y=39
        pixel_data[39][48] = 4'b1101; // x=48, y=39
        pixel_data[39][49] = 4'b0001; // x=49, y=39
        pixel_data[39][50] = 4'b0001; // x=50, y=39
        pixel_data[39][51] = 4'b0001; // x=51, y=39
        pixel_data[39][52] = 4'b1101; // x=52, y=39
        pixel_data[39][53] = 4'b1101; // x=53, y=39
        pixel_data[39][54] = 4'b1011; // x=54, y=39
        pixel_data[39][55] = 4'b1001; // x=55, y=39
        pixel_data[39][56] = 4'b0000; // x=56, y=39
        pixel_data[39][57] = 4'b0000; // x=57, y=39
        pixel_data[39][58] = 4'b0111; // x=58, y=39
        pixel_data[39][59] = 4'b0000; // x=59, y=39
        pixel_data[39][60] = 4'b0000; // x=60, y=39
        pixel_data[39][61] = 4'b0111; // x=61, y=39
        pixel_data[39][62] = 4'b0110; // x=62, y=39
        pixel_data[39][63] = 4'b1000; // x=63, y=39
        pixel_data[39][64] = 4'b1101; // x=64, y=39
        pixel_data[39][65] = 4'b1101; // x=65, y=39
        pixel_data[39][66] = 4'b1101; // x=66, y=39
        pixel_data[39][67] = 4'b0001; // x=67, y=39
        pixel_data[39][68] = 4'b0001; // x=68, y=39
        pixel_data[39][69] = 4'b0001; // x=69, y=39
        pixel_data[39][70] = 4'b1101; // x=70, y=39
        pixel_data[39][71] = 4'b1101; // x=71, y=39
        pixel_data[39][72] = 4'b1101; // x=72, y=39
        pixel_data[39][73] = 4'b0001; // x=73, y=39
        pixel_data[39][74] = 4'b0001; // x=74, y=39
        pixel_data[39][75] = 4'b1101; // x=75, y=39
        pixel_data[39][76] = 4'b1101; // x=76, y=39
        pixel_data[39][77] = 4'b1101; // x=77, y=39
        pixel_data[39][78] = 4'b0011; // x=78, y=39
        pixel_data[39][79] = 4'b0100; // x=79, y=39
        pixel_data[39][80] = 4'b0111; // x=80, y=39
        pixel_data[39][81] = 4'b0000; // x=81, y=39
        pixel_data[39][82] = 4'b0111; // x=82, y=39
        pixel_data[39][83] = 4'b0111; // x=83, y=39
        pixel_data[39][84] = 4'b0111; // x=84, y=39
        pixel_data[39][85] = 4'b0111; // x=85, y=39
        pixel_data[39][86] = 4'b0111; // x=86, y=39
        pixel_data[39][87] = 4'b0110; // x=87, y=39
        pixel_data[39][88] = 4'b1011; // x=88, y=39
        pixel_data[39][89] = 4'b0001; // x=89, y=39
        pixel_data[39][90] = 4'b0001; // x=90, y=39
        pixel_data[39][91] = 4'b0001; // x=91, y=39
        pixel_data[39][92] = 4'b0001; // x=92, y=39
        pixel_data[39][93] = 4'b1001; // x=93, y=39
        pixel_data[39][94] = 4'b0111; // x=94, y=39
        pixel_data[39][95] = 4'b0000; // x=95, y=39
        pixel_data[39][96] = 4'b0111; // x=96, y=39
        pixel_data[39][97] = 4'b0111; // x=97, y=39
        pixel_data[39][98] = 4'b0111; // x=98, y=39
        pixel_data[39][99] = 4'b0111; // x=99, y=39
        pixel_data[39][100] = 4'b0111; // x=100, y=39
        pixel_data[39][101] = 4'b0111; // x=101, y=39
        pixel_data[39][102] = 4'b0111; // x=102, y=39
        pixel_data[39][103] = 4'b0111; // x=103, y=39
        pixel_data[39][104] = 4'b0000; // x=104, y=39
        pixel_data[39][105] = 4'b0000; // x=105, y=39
        pixel_data[39][106] = 4'b0111; // x=106, y=39
        pixel_data[39][107] = 4'b1010; // x=107, y=39
        pixel_data[39][108] = 4'b1011; // x=108, y=39
        pixel_data[39][109] = 4'b1101; // x=109, y=39
        pixel_data[39][110] = 4'b1101; // x=110, y=39
        pixel_data[39][111] = 4'b1101; // x=111, y=39
        pixel_data[39][112] = 4'b0001; // x=112, y=39
        pixel_data[39][113] = 4'b0001; // x=113, y=39
        pixel_data[39][114] = 4'b1101; // x=114, y=39
        pixel_data[39][115] = 4'b1101; // x=115, y=39
        pixel_data[39][116] = 4'b1101; // x=116, y=39
        pixel_data[39][117] = 4'b1101; // x=117, y=39
        pixel_data[39][118] = 4'b0001; // x=118, y=39
        pixel_data[39][119] = 4'b0001; // x=119, y=39
        pixel_data[39][120] = 4'b0001; // x=120, y=39
        pixel_data[39][121] = 4'b1101; // x=121, y=39
        pixel_data[39][122] = 4'b1101; // x=122, y=39
        pixel_data[39][123] = 4'b0011; // x=123, y=39
        pixel_data[39][124] = 4'b0010; // x=124, y=39
        pixel_data[39][125] = 4'b0000; // x=125, y=39
        pixel_data[39][126] = 4'b0111; // x=126, y=39
        pixel_data[39][127] = 4'b0111; // x=127, y=39
        pixel_data[39][128] = 4'b0111; // x=128, y=39
        pixel_data[39][129] = 4'b0111; // x=129, y=39
        pixel_data[39][130] = 4'b0111; // x=130, y=39
        pixel_data[39][131] = 4'b0111; // x=131, y=39
        pixel_data[39][132] = 4'b0111; // x=132, y=39
        pixel_data[39][133] = 4'b0111; // x=133, y=39
        pixel_data[39][134] = 4'b0111; // x=134, y=39
        pixel_data[39][135] = 4'b0111; // x=135, y=39
        pixel_data[39][136] = 4'b0111; // x=136, y=39
        pixel_data[39][137] = 4'b0111; // x=137, y=39
        pixel_data[39][138] = 4'b0111; // x=138, y=39
        pixel_data[39][139] = 4'b0111; // x=139, y=39
        pixel_data[39][140] = 4'b0000; // x=140, y=39
        pixel_data[39][141] = 4'b0111; // x=141, y=39
        pixel_data[39][142] = 4'b0101; // x=142, y=39
        pixel_data[39][143] = 4'b1101; // x=143, y=39
        pixel_data[39][144] = 4'b0001; // x=144, y=39
        pixel_data[39][145] = 4'b1101; // x=145, y=39
        pixel_data[39][146] = 4'b0001; // x=146, y=39
        pixel_data[39][147] = 4'b1101; // x=147, y=39
        pixel_data[39][148] = 4'b0011; // x=148, y=39
        pixel_data[39][149] = 4'b0000; // x=149, y=39
        pixel_data[39][150] = 4'b0111; // x=150, y=39
        pixel_data[39][151] = 4'b0000; // x=151, y=39
        pixel_data[39][152] = 4'b0000; // x=152, y=39
        pixel_data[39][153] = 4'b0111; // x=153, y=39
        pixel_data[39][154] = 4'b0111; // x=154, y=39
        pixel_data[39][155] = 4'b0111; // x=155, y=39
        pixel_data[39][156] = 4'b0111; // x=156, y=39
        pixel_data[39][157] = 4'b0111; // x=157, y=39
        pixel_data[39][158] = 4'b0111; // x=158, y=39
        pixel_data[39][159] = 4'b0111; // x=159, y=39
        pixel_data[39][160] = 4'b0111; // x=160, y=39
        pixel_data[39][161] = 4'b0111; // x=161, y=39
        pixel_data[39][162] = 4'b0111; // x=162, y=39
        pixel_data[39][163] = 4'b0111; // x=163, y=39
        pixel_data[39][164] = 4'b0111; // x=164, y=39
        pixel_data[39][165] = 4'b0111; // x=165, y=39
        pixel_data[39][166] = 4'b0111; // x=166, y=39
        pixel_data[39][167] = 4'b0111; // x=167, y=39
        pixel_data[39][168] = 4'b0111; // x=168, y=39
        pixel_data[39][169] = 4'b0111; // x=169, y=39
        pixel_data[39][170] = 4'b0111; // x=170, y=39
        pixel_data[39][171] = 4'b0111; // x=171, y=39
        pixel_data[39][172] = 4'b0111; // x=172, y=39
        pixel_data[39][173] = 4'b0111; // x=173, y=39
        pixel_data[39][174] = 4'b0111; // x=174, y=39
        pixel_data[39][175] = 4'b0111; // x=175, y=39
        pixel_data[39][176] = 4'b0111; // x=176, y=39
        pixel_data[39][177] = 4'b0111; // x=177, y=39
        pixel_data[39][178] = 4'b0111; // x=178, y=39
        pixel_data[39][179] = 4'b0111; // x=179, y=39
        pixel_data[40][0] = 4'b0111; // x=0, y=40
        pixel_data[40][1] = 4'b0111; // x=1, y=40
        pixel_data[40][2] = 4'b0111; // x=2, y=40
        pixel_data[40][3] = 4'b0111; // x=3, y=40
        pixel_data[40][4] = 4'b0111; // x=4, y=40
        pixel_data[40][5] = 4'b0111; // x=5, y=40
        pixel_data[40][6] = 4'b0111; // x=6, y=40
        pixel_data[40][7] = 4'b0111; // x=7, y=40
        pixel_data[40][8] = 4'b0111; // x=8, y=40
        pixel_data[40][9] = 4'b0000; // x=9, y=40
        pixel_data[40][10] = 4'b0000; // x=10, y=40
        pixel_data[40][11] = 4'b0111; // x=11, y=40
        pixel_data[40][12] = 4'b0110; // x=12, y=40
        pixel_data[40][13] = 4'b0101; // x=13, y=40
        pixel_data[40][14] = 4'b0011; // x=14, y=40
        pixel_data[40][15] = 4'b1101; // x=15, y=40
        pixel_data[40][16] = 4'b1101; // x=16, y=40
        pixel_data[40][17] = 4'b1101; // x=17, y=40
        pixel_data[40][18] = 4'b1101; // x=18, y=40
        pixel_data[40][19] = 4'b1101; // x=19, y=40
        pixel_data[40][20] = 4'b1101; // x=20, y=40
        pixel_data[40][21] = 4'b1101; // x=21, y=40
        pixel_data[40][22] = 4'b1101; // x=22, y=40
        pixel_data[40][23] = 4'b1101; // x=23, y=40
        pixel_data[40][24] = 4'b1101; // x=24, y=40
        pixel_data[40][25] = 4'b0001; // x=25, y=40
        pixel_data[40][26] = 4'b0011; // x=26, y=40
        pixel_data[40][27] = 4'b1010; // x=27, y=40
        pixel_data[40][28] = 4'b1110; // x=28, y=40
        pixel_data[40][29] = 4'b0111; // x=29, y=40
        pixel_data[40][30] = 4'b0000; // x=30, y=40
        pixel_data[40][31] = 4'b0111; // x=31, y=40
        pixel_data[40][32] = 4'b0111; // x=32, y=40
        pixel_data[40][33] = 4'b0111; // x=33, y=40
        pixel_data[40][34] = 4'b0111; // x=34, y=40
        pixel_data[40][35] = 4'b0111; // x=35, y=40
        pixel_data[40][36] = 4'b0000; // x=36, y=40
        pixel_data[40][37] = 4'b0111; // x=37, y=40
        pixel_data[40][38] = 4'b0000; // x=38, y=40
        pixel_data[40][39] = 4'b0111; // x=39, y=40
        pixel_data[40][40] = 4'b0110; // x=40, y=40
        pixel_data[40][41] = 4'b0101; // x=41, y=40
        pixel_data[40][42] = 4'b1011; // x=42, y=40
        pixel_data[40][43] = 4'b1101; // x=43, y=40
        pixel_data[40][44] = 4'b1101; // x=44, y=40
        pixel_data[40][45] = 4'b1101; // x=45, y=40
        pixel_data[40][46] = 4'b1101; // x=46, y=40
        pixel_data[40][47] = 4'b1101; // x=47, y=40
        pixel_data[40][48] = 4'b1101; // x=48, y=40
        pixel_data[40][49] = 4'b1101; // x=49, y=40
        pixel_data[40][50] = 4'b1101; // x=50, y=40
        pixel_data[40][51] = 4'b1101; // x=51, y=40
        pixel_data[40][52] = 4'b0011; // x=52, y=40
        pixel_data[40][53] = 4'b0010; // x=53, y=40
        pixel_data[40][54] = 4'b1110; // x=54, y=40
        pixel_data[40][55] = 4'b0111; // x=55, y=40
        pixel_data[40][56] = 4'b0000; // x=56, y=40
        pixel_data[40][57] = 4'b0000; // x=57, y=40
        pixel_data[40][58] = 4'b0000; // x=58, y=40
        pixel_data[40][59] = 4'b0000; // x=59, y=40
        pixel_data[40][60] = 4'b0111; // x=60, y=40
        pixel_data[40][61] = 4'b0000; // x=61, y=40
        pixel_data[40][62] = 4'b0111; // x=62, y=40
        pixel_data[40][63] = 4'b0111; // x=63, y=40
        pixel_data[40][64] = 4'b1001; // x=64, y=40
        pixel_data[40][65] = 4'b1100; // x=65, y=40
        pixel_data[40][66] = 4'b0001; // x=66, y=40
        pixel_data[40][67] = 4'b1101; // x=67, y=40
        pixel_data[40][68] = 4'b1101; // x=68, y=40
        pixel_data[40][69] = 4'b1101; // x=69, y=40
        pixel_data[40][70] = 4'b1101; // x=70, y=40
        pixel_data[40][71] = 4'b1101; // x=71, y=40
        pixel_data[40][72] = 4'b1101; // x=72, y=40
        pixel_data[40][73] = 4'b1101; // x=73, y=40
        pixel_data[40][74] = 4'b1101; // x=74, y=40
        pixel_data[40][75] = 4'b0001; // x=75, y=40
        pixel_data[40][76] = 4'b0011; // x=76, y=40
        pixel_data[40][77] = 4'b1010; // x=77, y=40
        pixel_data[40][78] = 4'b0000; // x=78, y=40
        pixel_data[40][79] = 4'b0111; // x=79, y=40
        pixel_data[40][80] = 4'b0000; // x=80, y=40
        pixel_data[40][81] = 4'b0111; // x=81, y=40
        pixel_data[40][82] = 4'b0111; // x=82, y=40
        pixel_data[40][83] = 4'b0111; // x=83, y=40
        pixel_data[40][84] = 4'b0111; // x=84, y=40
        pixel_data[40][85] = 4'b0111; // x=85, y=40
        pixel_data[40][86] = 4'b0111; // x=86, y=40
        pixel_data[40][87] = 4'b0110; // x=87, y=40
        pixel_data[40][88] = 4'b1101; // x=88, y=40
        pixel_data[40][89] = 4'b1101; // x=89, y=40
        pixel_data[40][90] = 4'b1101; // x=90, y=40
        pixel_data[40][91] = 4'b1101; // x=91, y=40
        pixel_data[40][92] = 4'b1101; // x=92, y=40
        pixel_data[40][93] = 4'b1010; // x=93, y=40
        pixel_data[40][94] = 4'b0111; // x=94, y=40
        pixel_data[40][95] = 4'b0000; // x=95, y=40
        pixel_data[40][96] = 4'b0111; // x=96, y=40
        pixel_data[40][97] = 4'b0111; // x=97, y=40
        pixel_data[40][98] = 4'b0111; // x=98, y=40
        pixel_data[40][99] = 4'b0111; // x=99, y=40
        pixel_data[40][100] = 4'b0111; // x=100, y=40
        pixel_data[40][101] = 4'b0111; // x=101, y=40
        pixel_data[40][102] = 4'b0111; // x=102, y=40
        pixel_data[40][103] = 4'b0111; // x=103, y=40
        pixel_data[40][104] = 4'b0000; // x=104, y=40
        pixel_data[40][105] = 4'b0000; // x=105, y=40
        pixel_data[40][106] = 4'b0000; // x=106, y=40
        pixel_data[40][107] = 4'b0111; // x=107, y=40
        pixel_data[40][108] = 4'b1110; // x=108, y=40
        pixel_data[40][109] = 4'b0010; // x=109, y=40
        pixel_data[40][110] = 4'b0011; // x=110, y=40
        pixel_data[40][111] = 4'b1101; // x=111, y=40
        pixel_data[40][112] = 4'b1101; // x=112, y=40
        pixel_data[40][113] = 4'b1101; // x=113, y=40
        pixel_data[40][114] = 4'b1101; // x=114, y=40
        pixel_data[40][115] = 4'b1101; // x=115, y=40
        pixel_data[40][116] = 4'b1101; // x=116, y=40
        pixel_data[40][117] = 4'b1101; // x=117, y=40
        pixel_data[40][118] = 4'b1101; // x=118, y=40
        pixel_data[40][119] = 4'b1101; // x=119, y=40
        pixel_data[40][120] = 4'b0001; // x=120, y=40
        pixel_data[40][121] = 4'b1100; // x=121, y=40
        pixel_data[40][122] = 4'b0010; // x=122, y=40
        pixel_data[40][123] = 4'b1110; // x=123, y=40
        pixel_data[40][124] = 4'b0111; // x=124, y=40
        pixel_data[40][125] = 4'b0000; // x=125, y=40
        pixel_data[40][126] = 4'b0111; // x=126, y=40
        pixel_data[40][127] = 4'b0111; // x=127, y=40
        pixel_data[40][128] = 4'b0111; // x=128, y=40
        pixel_data[40][129] = 4'b0111; // x=129, y=40
        pixel_data[40][130] = 4'b0111; // x=130, y=40
        pixel_data[40][131] = 4'b0111; // x=131, y=40
        pixel_data[40][132] = 4'b0111; // x=132, y=40
        pixel_data[40][133] = 4'b0111; // x=133, y=40
        pixel_data[40][134] = 4'b0111; // x=134, y=40
        pixel_data[40][135] = 4'b0111; // x=135, y=40
        pixel_data[40][136] = 4'b0111; // x=136, y=40
        pixel_data[40][137] = 4'b0111; // x=137, y=40
        pixel_data[40][138] = 4'b0111; // x=138, y=40
        pixel_data[40][139] = 4'b0111; // x=139, y=40
        pixel_data[40][140] = 4'b0000; // x=140, y=40
        pixel_data[40][141] = 4'b0111; // x=141, y=40
        pixel_data[40][142] = 4'b0100; // x=142, y=40
        pixel_data[40][143] = 4'b0001; // x=143, y=40
        pixel_data[40][144] = 4'b1101; // x=144, y=40
        pixel_data[40][145] = 4'b1101; // x=145, y=40
        pixel_data[40][146] = 4'b1101; // x=146, y=40
        pixel_data[40][147] = 4'b1101; // x=147, y=40
        pixel_data[40][148] = 4'b1010; // x=148, y=40
        pixel_data[40][149] = 4'b0111; // x=149, y=40
        pixel_data[40][150] = 4'b0000; // x=150, y=40
        pixel_data[40][151] = 4'b0111; // x=151, y=40
        pixel_data[40][152] = 4'b0111; // x=152, y=40
        pixel_data[40][153] = 4'b0111; // x=153, y=40
        pixel_data[40][154] = 4'b0111; // x=154, y=40
        pixel_data[40][155] = 4'b0111; // x=155, y=40
        pixel_data[40][156] = 4'b0111; // x=156, y=40
        pixel_data[40][157] = 4'b0111; // x=157, y=40
        pixel_data[40][158] = 4'b0111; // x=158, y=40
        pixel_data[40][159] = 4'b0111; // x=159, y=40
        pixel_data[40][160] = 4'b0111; // x=160, y=40
        pixel_data[40][161] = 4'b0111; // x=161, y=40
        pixel_data[40][162] = 4'b0111; // x=162, y=40
        pixel_data[40][163] = 4'b0111; // x=163, y=40
        pixel_data[40][164] = 4'b0111; // x=164, y=40
        pixel_data[40][165] = 4'b0111; // x=165, y=40
        pixel_data[40][166] = 4'b0111; // x=166, y=40
        pixel_data[40][167] = 4'b0111; // x=167, y=40
        pixel_data[40][168] = 4'b0111; // x=168, y=40
        pixel_data[40][169] = 4'b0111; // x=169, y=40
        pixel_data[40][170] = 4'b0111; // x=170, y=40
        pixel_data[40][171] = 4'b0111; // x=171, y=40
        pixel_data[40][172] = 4'b0111; // x=172, y=40
        pixel_data[40][173] = 4'b0111; // x=173, y=40
        pixel_data[40][174] = 4'b0111; // x=174, y=40
        pixel_data[40][175] = 4'b0111; // x=175, y=40
        pixel_data[40][176] = 4'b0111; // x=176, y=40
        pixel_data[40][177] = 4'b0111; // x=177, y=40
        pixel_data[40][178] = 4'b0111; // x=178, y=40
        pixel_data[40][179] = 4'b0111; // x=179, y=40
        pixel_data[41][0] = 4'b0111; // x=0, y=41
        pixel_data[41][1] = 4'b0111; // x=1, y=41
        pixel_data[41][2] = 4'b0111; // x=2, y=41
        pixel_data[41][3] = 4'b0111; // x=3, y=41
        pixel_data[41][4] = 4'b0111; // x=4, y=41
        pixel_data[41][5] = 4'b0111; // x=5, y=41
        pixel_data[41][6] = 4'b0111; // x=6, y=41
        pixel_data[41][7] = 4'b0111; // x=7, y=41
        pixel_data[41][8] = 4'b0111; // x=8, y=41
        pixel_data[41][9] = 4'b0000; // x=9, y=41
        pixel_data[41][10] = 4'b0000; // x=10, y=41
        pixel_data[41][11] = 4'b0000; // x=11, y=41
        pixel_data[41][12] = 4'b0111; // x=12, y=41
        pixel_data[41][13] = 4'b0111; // x=13, y=41
        pixel_data[41][14] = 4'b0000; // x=14, y=41
        pixel_data[41][15] = 4'b0100; // x=15, y=41
        pixel_data[41][16] = 4'b1010; // x=16, y=41
        pixel_data[41][17] = 4'b0101; // x=17, y=41
        pixel_data[41][18] = 4'b1000; // x=18, y=41
        pixel_data[41][19] = 4'b1100; // x=19, y=41
        pixel_data[41][20] = 4'b1100; // x=20, y=41
        pixel_data[41][21] = 4'b1000; // x=21, y=41
        pixel_data[41][22] = 4'b1111; // x=22, y=41
        pixel_data[41][23] = 4'b0101; // x=23, y=41
        pixel_data[41][24] = 4'b1010; // x=24, y=41
        pixel_data[41][25] = 4'b0110; // x=25, y=41
        pixel_data[41][26] = 4'b0000; // x=26, y=41
        pixel_data[41][27] = 4'b0111; // x=27, y=41
        pixel_data[41][28] = 4'b0111; // x=28, y=41
        pixel_data[41][29] = 4'b0000; // x=29, y=41
        pixel_data[41][30] = 4'b0000; // x=30, y=41
        pixel_data[41][31] = 4'b0000; // x=31, y=41
        pixel_data[41][32] = 4'b0111; // x=32, y=41
        pixel_data[41][33] = 4'b0111; // x=33, y=41
        pixel_data[41][34] = 4'b0111; // x=34, y=41
        pixel_data[41][35] = 4'b0111; // x=35, y=41
        pixel_data[41][36] = 4'b0111; // x=36, y=41
        pixel_data[41][37] = 4'b0000; // x=37, y=41
        pixel_data[41][38] = 4'b0000; // x=38, y=41
        pixel_data[41][39] = 4'b0000; // x=39, y=41
        pixel_data[41][40] = 4'b0111; // x=40, y=41
        pixel_data[41][41] = 4'b0111; // x=41, y=41
        pixel_data[41][42] = 4'b1110; // x=42, y=41
        pixel_data[41][43] = 4'b1001; // x=43, y=41
        pixel_data[41][44] = 4'b0101; // x=44, y=41
        pixel_data[41][45] = 4'b1111; // x=45, y=41
        pixel_data[41][46] = 4'b1100; // x=46, y=41
        pixel_data[41][47] = 4'b1100; // x=47, y=41
        pixel_data[41][48] = 4'b1000; // x=48, y=41
        pixel_data[41][49] = 4'b0101; // x=49, y=41
        pixel_data[41][50] = 4'b0010; // x=50, y=41
        pixel_data[41][51] = 4'b0100; // x=51, y=41
        pixel_data[41][52] = 4'b0000; // x=52, y=41
        pixel_data[41][53] = 4'b0111; // x=53, y=41
        pixel_data[41][54] = 4'b0111; // x=54, y=41
        pixel_data[41][55] = 4'b0000; // x=55, y=41
        pixel_data[41][56] = 4'b0000; // x=56, y=41
        pixel_data[41][57] = 4'b0111; // x=57, y=41
        pixel_data[41][58] = 4'b0111; // x=58, y=41
        pixel_data[41][59] = 4'b0000; // x=59, y=41
        pixel_data[41][60] = 4'b0111; // x=60, y=41
        pixel_data[41][61] = 4'b0000; // x=61, y=41
        pixel_data[41][62] = 4'b0000; // x=62, y=41
        pixel_data[41][63] = 4'b0000; // x=63, y=41
        pixel_data[41][64] = 4'b0111; // x=64, y=41
        pixel_data[41][65] = 4'b0111; // x=65, y=41
        pixel_data[41][66] = 4'b0110; // x=66, y=41
        pixel_data[41][67] = 4'b1010; // x=67, y=41
        pixel_data[41][68] = 4'b0101; // x=68, y=41
        pixel_data[41][69] = 4'b1111; // x=69, y=41
        pixel_data[41][70] = 4'b1100; // x=70, y=41
        pixel_data[41][71] = 4'b1100; // x=71, y=41
        pixel_data[41][72] = 4'b1000; // x=72, y=41
        pixel_data[41][73] = 4'b0101; // x=73, y=41
        pixel_data[41][74] = 4'b0010; // x=74, y=41
        pixel_data[41][75] = 4'b0100; // x=75, y=41
        pixel_data[41][76] = 4'b0000; // x=76, y=41
        pixel_data[41][77] = 4'b0111; // x=77, y=41
        pixel_data[41][78] = 4'b0111; // x=78, y=41
        pixel_data[41][79] = 4'b0000; // x=79, y=41
        pixel_data[41][80] = 4'b0111; // x=80, y=41
        pixel_data[41][81] = 4'b0111; // x=81, y=41
        pixel_data[41][82] = 4'b0111; // x=82, y=41
        pixel_data[41][83] = 4'b0111; // x=83, y=41
        pixel_data[41][84] = 4'b0111; // x=84, y=41
        pixel_data[41][85] = 4'b0111; // x=85, y=41
        pixel_data[41][86] = 4'b0000; // x=86, y=41
        pixel_data[41][87] = 4'b1110; // x=87, y=41
        pixel_data[41][88] = 4'b0010; // x=88, y=41
        pixel_data[41][89] = 4'b0010; // x=89, y=41
        pixel_data[41][90] = 4'b0010; // x=90, y=41
        pixel_data[41][91] = 4'b0010; // x=91, y=41
        pixel_data[41][92] = 4'b0010; // x=92, y=41
        pixel_data[41][93] = 4'b0110; // x=93, y=41
        pixel_data[41][94] = 4'b0111; // x=94, y=41
        pixel_data[41][95] = 4'b0111; // x=95, y=41
        pixel_data[41][96] = 4'b0111; // x=96, y=41
        pixel_data[41][97] = 4'b0111; // x=97, y=41
        pixel_data[41][98] = 4'b0111; // x=98, y=41
        pixel_data[41][99] = 4'b0111; // x=99, y=41
        pixel_data[41][100] = 4'b0111; // x=100, y=41
        pixel_data[41][101] = 4'b0111; // x=101, y=41
        pixel_data[41][102] = 4'b0111; // x=102, y=41
        pixel_data[41][103] = 4'b0111; // x=103, y=41
        pixel_data[41][104] = 4'b0000; // x=104, y=41
        pixel_data[41][105] = 4'b0000; // x=105, y=41
        pixel_data[41][106] = 4'b0111; // x=106, y=41
        pixel_data[41][107] = 4'b0000; // x=107, y=41
        pixel_data[41][108] = 4'b0111; // x=108, y=41
        pixel_data[41][109] = 4'b0111; // x=109, y=41
        pixel_data[41][110] = 4'b0000; // x=110, y=41
        pixel_data[41][111] = 4'b0100; // x=111, y=41
        pixel_data[41][112] = 4'b0010; // x=112, y=41
        pixel_data[41][113] = 4'b0101; // x=113, y=41
        pixel_data[41][114] = 4'b1111; // x=114, y=41
        pixel_data[41][115] = 4'b1100; // x=115, y=41
        pixel_data[41][116] = 4'b1100; // x=116, y=41
        pixel_data[41][117] = 4'b1111; // x=117, y=41
        pixel_data[41][118] = 4'b0101; // x=118, y=41
        pixel_data[41][119] = 4'b1010; // x=119, y=41
        pixel_data[41][120] = 4'b0110; // x=120, y=41
        pixel_data[41][121] = 4'b0000; // x=121, y=41
        pixel_data[41][122] = 4'b0111; // x=122, y=41
        pixel_data[41][123] = 4'b0111; // x=123, y=41
        pixel_data[41][124] = 4'b0000; // x=124, y=41
        pixel_data[41][125] = 4'b0000; // x=125, y=41
        pixel_data[41][126] = 4'b0111; // x=126, y=41
        pixel_data[41][127] = 4'b0111; // x=127, y=41
        pixel_data[41][128] = 4'b0111; // x=128, y=41
        pixel_data[41][129] = 4'b0111; // x=129, y=41
        pixel_data[41][130] = 4'b0111; // x=130, y=41
        pixel_data[41][131] = 4'b0111; // x=131, y=41
        pixel_data[41][132] = 4'b0111; // x=132, y=41
        pixel_data[41][133] = 4'b0111; // x=133, y=41
        pixel_data[41][134] = 4'b0111; // x=134, y=41
        pixel_data[41][135] = 4'b0111; // x=135, y=41
        pixel_data[41][136] = 4'b0111; // x=136, y=41
        pixel_data[41][137] = 4'b0111; // x=137, y=41
        pixel_data[41][138] = 4'b0111; // x=138, y=41
        pixel_data[41][139] = 4'b0111; // x=139, y=41
        pixel_data[41][140] = 4'b0111; // x=140, y=41
        pixel_data[41][141] = 4'b0111; // x=141, y=41
        pixel_data[41][142] = 4'b0111; // x=142, y=41
        pixel_data[41][143] = 4'b0100; // x=143, y=41
        pixel_data[41][144] = 4'b1111; // x=144, y=41
        pixel_data[41][145] = 4'b1100; // x=145, y=41
        pixel_data[41][146] = 4'b1000; // x=146, y=41
        pixel_data[41][147] = 4'b1001; // x=147, y=41
        pixel_data[41][148] = 4'b0111; // x=148, y=41
        pixel_data[41][149] = 4'b0000; // x=149, y=41
        pixel_data[41][150] = 4'b0111; // x=150, y=41
        pixel_data[41][151] = 4'b0111; // x=151, y=41
        pixel_data[41][152] = 4'b0111; // x=152, y=41
        pixel_data[41][153] = 4'b0111; // x=153, y=41
        pixel_data[41][154] = 4'b0111; // x=154, y=41
        pixel_data[41][155] = 4'b0111; // x=155, y=41
        pixel_data[41][156] = 4'b0111; // x=156, y=41
        pixel_data[41][157] = 4'b0111; // x=157, y=41
        pixel_data[41][158] = 4'b0111; // x=158, y=41
        pixel_data[41][159] = 4'b0111; // x=159, y=41
        pixel_data[41][160] = 4'b0111; // x=160, y=41
        pixel_data[41][161] = 4'b0111; // x=161, y=41
        pixel_data[41][162] = 4'b0111; // x=162, y=41
        pixel_data[41][163] = 4'b0111; // x=163, y=41
        pixel_data[41][164] = 4'b0111; // x=164, y=41
        pixel_data[41][165] = 4'b0111; // x=165, y=41
        pixel_data[41][166] = 4'b0111; // x=166, y=41
        pixel_data[41][167] = 4'b0111; // x=167, y=41
        pixel_data[41][168] = 4'b0111; // x=168, y=41
        pixel_data[41][169] = 4'b0111; // x=169, y=41
        pixel_data[41][170] = 4'b0111; // x=170, y=41
        pixel_data[41][171] = 4'b0111; // x=171, y=41
        pixel_data[41][172] = 4'b0111; // x=172, y=41
        pixel_data[41][173] = 4'b0111; // x=173, y=41
        pixel_data[41][174] = 4'b0111; // x=174, y=41
        pixel_data[41][175] = 4'b0111; // x=175, y=41
        pixel_data[41][176] = 4'b0111; // x=176, y=41
        pixel_data[41][177] = 4'b0111; // x=177, y=41
        pixel_data[41][178] = 4'b0111; // x=178, y=41
        pixel_data[41][179] = 4'b0111; // x=179, y=41
        pixel_data[42][0] = 4'b0111; // x=0, y=42
        pixel_data[42][1] = 4'b0111; // x=1, y=42
        pixel_data[42][2] = 4'b0111; // x=2, y=42
        pixel_data[42][3] = 4'b0111; // x=3, y=42
        pixel_data[42][4] = 4'b0111; // x=4, y=42
        pixel_data[42][5] = 4'b0111; // x=5, y=42
        pixel_data[42][6] = 4'b0111; // x=6, y=42
        pixel_data[42][7] = 4'b0111; // x=7, y=42
        pixel_data[42][8] = 4'b0111; // x=8, y=42
        pixel_data[42][9] = 4'b0111; // x=9, y=42
        pixel_data[42][10] = 4'b0111; // x=10, y=42
        pixel_data[42][11] = 4'b0000; // x=11, y=42
        pixel_data[42][12] = 4'b0000; // x=12, y=42
        pixel_data[42][13] = 4'b0000; // x=13, y=42
        pixel_data[42][14] = 4'b0111; // x=14, y=42
        pixel_data[42][15] = 4'b0111; // x=15, y=42
        pixel_data[42][16] = 4'b0111; // x=16, y=42
        pixel_data[42][17] = 4'b0111; // x=17, y=42
        pixel_data[42][18] = 4'b0111; // x=18, y=42
        pixel_data[42][19] = 4'b0111; // x=19, y=42
        pixel_data[42][20] = 4'b0111; // x=20, y=42
        pixel_data[42][21] = 4'b0111; // x=21, y=42
        pixel_data[42][22] = 4'b0111; // x=22, y=42
        pixel_data[42][23] = 4'b0111; // x=23, y=42
        pixel_data[42][24] = 4'b0111; // x=24, y=42
        pixel_data[42][25] = 4'b0111; // x=25, y=42
        pixel_data[42][26] = 4'b0111; // x=26, y=42
        pixel_data[42][27] = 4'b0000; // x=27, y=42
        pixel_data[42][28] = 4'b0111; // x=28, y=42
        pixel_data[42][29] = 4'b0111; // x=29, y=42
        pixel_data[42][30] = 4'b0111; // x=30, y=42
        pixel_data[42][31] = 4'b0111; // x=31, y=42
        pixel_data[42][32] = 4'b0111; // x=32, y=42
        pixel_data[42][33] = 4'b0111; // x=33, y=42
        pixel_data[42][34] = 4'b0111; // x=34, y=42
        pixel_data[42][35] = 4'b0111; // x=35, y=42
        pixel_data[42][36] = 4'b0111; // x=36, y=42
        pixel_data[42][37] = 4'b0111; // x=37, y=42
        pixel_data[42][38] = 4'b0000; // x=38, y=42
        pixel_data[42][39] = 4'b0111; // x=39, y=42
        pixel_data[42][40] = 4'b0000; // x=40, y=42
        pixel_data[42][41] = 4'b0000; // x=41, y=42
        pixel_data[42][42] = 4'b0111; // x=42, y=42
        pixel_data[42][43] = 4'b0111; // x=43, y=42
        pixel_data[42][44] = 4'b0111; // x=44, y=42
        pixel_data[42][45] = 4'b0111; // x=45, y=42
        pixel_data[42][46] = 4'b0111; // x=46, y=42
        pixel_data[42][47] = 4'b0111; // x=47, y=42
        pixel_data[42][48] = 4'b0111; // x=48, y=42
        pixel_data[42][49] = 4'b0111; // x=49, y=42
        pixel_data[42][50] = 4'b0111; // x=50, y=42
        pixel_data[42][51] = 4'b0111; // x=51, y=42
        pixel_data[42][52] = 4'b0111; // x=52, y=42
        pixel_data[42][53] = 4'b0000; // x=53, y=42
        pixel_data[42][54] = 4'b0000; // x=54, y=42
        pixel_data[42][55] = 4'b0111; // x=55, y=42
        pixel_data[42][56] = 4'b0111; // x=56, y=42
        pixel_data[42][57] = 4'b0111; // x=57, y=42
        pixel_data[42][58] = 4'b0111; // x=58, y=42
        pixel_data[42][59] = 4'b0111; // x=59, y=42
        pixel_data[42][60] = 4'b0111; // x=60, y=42
        pixel_data[42][61] = 4'b0111; // x=61, y=42
        pixel_data[42][62] = 4'b0111; // x=62, y=42
        pixel_data[42][63] = 4'b0111; // x=63, y=42
        pixel_data[42][64] = 4'b0000; // x=64, y=42
        pixel_data[42][65] = 4'b0111; // x=65, y=42
        pixel_data[42][66] = 4'b0111; // x=66, y=42
        pixel_data[42][67] = 4'b0111; // x=67, y=42
        pixel_data[42][68] = 4'b0111; // x=68, y=42
        pixel_data[42][69] = 4'b0111; // x=69, y=42
        pixel_data[42][70] = 4'b0111; // x=70, y=42
        pixel_data[42][71] = 4'b0111; // x=71, y=42
        pixel_data[42][72] = 4'b0111; // x=72, y=42
        pixel_data[42][73] = 4'b0111; // x=73, y=42
        pixel_data[42][74] = 4'b0111; // x=74, y=42
        pixel_data[42][75] = 4'b0111; // x=75, y=42
        pixel_data[42][76] = 4'b0111; // x=76, y=42
        pixel_data[42][77] = 4'b0000; // x=77, y=42
        pixel_data[42][78] = 4'b0111; // x=78, y=42
        pixel_data[42][79] = 4'b0111; // x=79, y=42
        pixel_data[42][80] = 4'b0111; // x=80, y=42
        pixel_data[42][81] = 4'b0111; // x=81, y=42
        pixel_data[42][82] = 4'b0111; // x=82, y=42
        pixel_data[42][83] = 4'b0111; // x=83, y=42
        pixel_data[42][84] = 4'b0111; // x=84, y=42
        pixel_data[42][85] = 4'b0111; // x=85, y=42
        pixel_data[42][86] = 4'b0111; // x=86, y=42
        pixel_data[42][87] = 4'b0111; // x=87, y=42
        pixel_data[42][88] = 4'b0111; // x=88, y=42
        pixel_data[42][89] = 4'b0111; // x=89, y=42
        pixel_data[42][90] = 4'b0111; // x=90, y=42
        pixel_data[42][91] = 4'b0111; // x=91, y=42
        pixel_data[42][92] = 4'b0111; // x=92, y=42
        pixel_data[42][93] = 4'b0111; // x=93, y=42
        pixel_data[42][94] = 4'b0111; // x=94, y=42
        pixel_data[42][95] = 4'b0111; // x=95, y=42
        pixel_data[42][96] = 4'b0111; // x=96, y=42
        pixel_data[42][97] = 4'b0111; // x=97, y=42
        pixel_data[42][98] = 4'b0111; // x=98, y=42
        pixel_data[42][99] = 4'b0111; // x=99, y=42
        pixel_data[42][100] = 4'b0111; // x=100, y=42
        pixel_data[42][101] = 4'b0111; // x=101, y=42
        pixel_data[42][102] = 4'b0111; // x=102, y=42
        pixel_data[42][103] = 4'b0111; // x=103, y=42
        pixel_data[42][104] = 4'b0111; // x=104, y=42
        pixel_data[42][105] = 4'b0111; // x=105, y=42
        pixel_data[42][106] = 4'b0111; // x=106, y=42
        pixel_data[42][107] = 4'b0111; // x=107, y=42
        pixel_data[42][108] = 4'b0111; // x=108, y=42
        pixel_data[42][109] = 4'b0000; // x=109, y=42
        pixel_data[42][110] = 4'b0111; // x=110, y=42
        pixel_data[42][111] = 4'b0111; // x=111, y=42
        pixel_data[42][112] = 4'b0111; // x=112, y=42
        pixel_data[42][113] = 4'b0111; // x=113, y=42
        pixel_data[42][114] = 4'b0111; // x=114, y=42
        pixel_data[42][115] = 4'b0111; // x=115, y=42
        pixel_data[42][116] = 4'b0111; // x=116, y=42
        pixel_data[42][117] = 4'b0111; // x=117, y=42
        pixel_data[42][118] = 4'b0111; // x=118, y=42
        pixel_data[42][119] = 4'b0111; // x=119, y=42
        pixel_data[42][120] = 4'b0111; // x=120, y=42
        pixel_data[42][121] = 4'b0111; // x=121, y=42
        pixel_data[42][122] = 4'b0000; // x=122, y=42
        pixel_data[42][123] = 4'b0111; // x=123, y=42
        pixel_data[42][124] = 4'b0111; // x=124, y=42
        pixel_data[42][125] = 4'b0111; // x=125, y=42
        pixel_data[42][126] = 4'b0111; // x=126, y=42
        pixel_data[42][127] = 4'b0111; // x=127, y=42
        pixel_data[42][128] = 4'b0111; // x=128, y=42
        pixel_data[42][129] = 4'b0111; // x=129, y=42
        pixel_data[42][130] = 4'b0111; // x=130, y=42
        pixel_data[42][131] = 4'b0111; // x=131, y=42
        pixel_data[42][132] = 4'b0111; // x=132, y=42
        pixel_data[42][133] = 4'b0111; // x=133, y=42
        pixel_data[42][134] = 4'b0111; // x=134, y=42
        pixel_data[42][135] = 4'b0111; // x=135, y=42
        pixel_data[42][136] = 4'b0111; // x=136, y=42
        pixel_data[42][137] = 4'b0111; // x=137, y=42
        pixel_data[42][138] = 4'b0111; // x=138, y=42
        pixel_data[42][139] = 4'b0111; // x=139, y=42
        pixel_data[42][140] = 4'b0111; // x=140, y=42
        pixel_data[42][141] = 4'b0111; // x=141, y=42
        pixel_data[42][142] = 4'b0000; // x=142, y=42
        pixel_data[42][143] = 4'b0111; // x=143, y=42
        pixel_data[42][144] = 4'b0111; // x=144, y=42
        pixel_data[42][145] = 4'b0111; // x=145, y=42
        pixel_data[42][146] = 4'b0111; // x=146, y=42
        pixel_data[42][147] = 4'b0111; // x=147, y=42
        pixel_data[42][148] = 4'b0111; // x=148, y=42
        pixel_data[42][149] = 4'b0111; // x=149, y=42
        pixel_data[42][150] = 4'b0111; // x=150, y=42
        pixel_data[42][151] = 4'b0111; // x=151, y=42
        pixel_data[42][152] = 4'b0111; // x=152, y=42
        pixel_data[42][153] = 4'b0111; // x=153, y=42
        pixel_data[42][154] = 4'b0111; // x=154, y=42
        pixel_data[42][155] = 4'b0111; // x=155, y=42
        pixel_data[42][156] = 4'b0111; // x=156, y=42
        pixel_data[42][157] = 4'b0111; // x=157, y=42
        pixel_data[42][158] = 4'b0111; // x=158, y=42
        pixel_data[42][159] = 4'b0111; // x=159, y=42
        pixel_data[42][160] = 4'b0111; // x=160, y=42
        pixel_data[42][161] = 4'b0111; // x=161, y=42
        pixel_data[42][162] = 4'b0111; // x=162, y=42
        pixel_data[42][163] = 4'b0111; // x=163, y=42
        pixel_data[42][164] = 4'b0111; // x=164, y=42
        pixel_data[42][165] = 4'b0111; // x=165, y=42
        pixel_data[42][166] = 4'b0111; // x=166, y=42
        pixel_data[42][167] = 4'b0111; // x=167, y=42
        pixel_data[42][168] = 4'b0111; // x=168, y=42
        pixel_data[42][169] = 4'b0111; // x=169, y=42
        pixel_data[42][170] = 4'b0111; // x=170, y=42
        pixel_data[42][171] = 4'b0111; // x=171, y=42
        pixel_data[42][172] = 4'b0111; // x=172, y=42
        pixel_data[42][173] = 4'b0111; // x=173, y=42
        pixel_data[42][174] = 4'b0111; // x=174, y=42
        pixel_data[42][175] = 4'b0111; // x=175, y=42
        pixel_data[42][176] = 4'b0111; // x=176, y=42
        pixel_data[42][177] = 4'b0111; // x=177, y=42
        pixel_data[42][178] = 4'b0111; // x=178, y=42
        pixel_data[42][179] = 4'b0111; // x=179, y=42
        pixel_data[43][0] = 4'b0111; // x=0, y=43
        pixel_data[43][1] = 4'b0111; // x=1, y=43
        pixel_data[43][2] = 4'b0111; // x=2, y=43
        pixel_data[43][3] = 4'b0111; // x=3, y=43
        pixel_data[43][4] = 4'b0111; // x=4, y=43
        pixel_data[43][5] = 4'b0111; // x=5, y=43
        pixel_data[43][6] = 4'b0111; // x=6, y=43
        pixel_data[43][7] = 4'b0111; // x=7, y=43
        pixel_data[43][8] = 4'b0111; // x=8, y=43
        pixel_data[43][9] = 4'b0111; // x=9, y=43
        pixel_data[43][10] = 4'b0111; // x=10, y=43
        pixel_data[43][11] = 4'b0111; // x=11, y=43
        pixel_data[43][12] = 4'b0111; // x=12, y=43
        pixel_data[43][13] = 4'b0111; // x=13, y=43
        pixel_data[43][14] = 4'b0111; // x=14, y=43
        pixel_data[43][15] = 4'b0111; // x=15, y=43
        pixel_data[43][16] = 4'b0000; // x=16, y=43
        pixel_data[43][17] = 4'b0000; // x=17, y=43
        pixel_data[43][18] = 4'b0111; // x=18, y=43
        pixel_data[43][19] = 4'b0111; // x=19, y=43
        pixel_data[43][20] = 4'b0111; // x=20, y=43
        pixel_data[43][21] = 4'b0111; // x=21, y=43
        pixel_data[43][22] = 4'b0111; // x=22, y=43
        pixel_data[43][23] = 4'b0000; // x=23, y=43
        pixel_data[43][24] = 4'b0000; // x=24, y=43
        pixel_data[43][25] = 4'b0111; // x=25, y=43
        pixel_data[43][26] = 4'b0111; // x=26, y=43
        pixel_data[43][27] = 4'b0111; // x=27, y=43
        pixel_data[43][28] = 4'b0111; // x=28, y=43
        pixel_data[43][29] = 4'b0111; // x=29, y=43
        pixel_data[43][30] = 4'b0111; // x=30, y=43
        pixel_data[43][31] = 4'b0111; // x=31, y=43
        pixel_data[43][32] = 4'b0111; // x=32, y=43
        pixel_data[43][33] = 4'b0111; // x=33, y=43
        pixel_data[43][34] = 4'b0111; // x=34, y=43
        pixel_data[43][35] = 4'b0111; // x=35, y=43
        pixel_data[43][36] = 4'b0111; // x=36, y=43
        pixel_data[43][37] = 4'b0111; // x=37, y=43
        pixel_data[43][38] = 4'b0111; // x=38, y=43
        pixel_data[43][39] = 4'b0111; // x=39, y=43
        pixel_data[43][40] = 4'b0111; // x=40, y=43
        pixel_data[43][41] = 4'b0111; // x=41, y=43
        pixel_data[43][42] = 4'b0111; // x=42, y=43
        pixel_data[43][43] = 4'b0000; // x=43, y=43
        pixel_data[43][44] = 4'b0000; // x=44, y=43
        pixel_data[43][45] = 4'b0111; // x=45, y=43
        pixel_data[43][46] = 4'b0111; // x=46, y=43
        pixel_data[43][47] = 4'b0111; // x=47, y=43
        pixel_data[43][48] = 4'b0111; // x=48, y=43
        pixel_data[43][49] = 4'b0000; // x=49, y=43
        pixel_data[43][50] = 4'b0000; // x=50, y=43
        pixel_data[43][51] = 4'b0111; // x=51, y=43
        pixel_data[43][52] = 4'b0111; // x=52, y=43
        pixel_data[43][53] = 4'b0111; // x=53, y=43
        pixel_data[43][54] = 4'b0111; // x=54, y=43
        pixel_data[43][55] = 4'b0111; // x=55, y=43
        pixel_data[43][56] = 4'b0111; // x=56, y=43
        pixel_data[43][57] = 4'b0111; // x=57, y=43
        pixel_data[43][58] = 4'b0111; // x=58, y=43
        pixel_data[43][59] = 4'b0111; // x=59, y=43
        pixel_data[43][60] = 4'b0111; // x=60, y=43
        pixel_data[43][61] = 4'b0111; // x=61, y=43
        pixel_data[43][62] = 4'b0111; // x=62, y=43
        pixel_data[43][63] = 4'b0111; // x=63, y=43
        pixel_data[43][64] = 4'b0111; // x=64, y=43
        pixel_data[43][65] = 4'b0111; // x=65, y=43
        pixel_data[43][66] = 4'b0111; // x=66, y=43
        pixel_data[43][67] = 4'b0000; // x=67, y=43
        pixel_data[43][68] = 4'b0000; // x=68, y=43
        pixel_data[43][69] = 4'b0111; // x=69, y=43
        pixel_data[43][70] = 4'b0111; // x=70, y=43
        pixel_data[43][71] = 4'b0111; // x=71, y=43
        pixel_data[43][72] = 4'b0111; // x=72, y=43
        pixel_data[43][73] = 4'b0000; // x=73, y=43
        pixel_data[43][74] = 4'b0000; // x=74, y=43
        pixel_data[43][75] = 4'b0111; // x=75, y=43
        pixel_data[43][76] = 4'b0111; // x=76, y=43
        pixel_data[43][77] = 4'b0111; // x=77, y=43
        pixel_data[43][78] = 4'b0111; // x=78, y=43
        pixel_data[43][79] = 4'b0111; // x=79, y=43
        pixel_data[43][80] = 4'b0111; // x=80, y=43
        pixel_data[43][81] = 4'b0111; // x=81, y=43
        pixel_data[43][82] = 4'b0111; // x=82, y=43
        pixel_data[43][83] = 4'b0111; // x=83, y=43
        pixel_data[43][84] = 4'b0111; // x=84, y=43
        pixel_data[43][85] = 4'b0111; // x=85, y=43
        pixel_data[43][86] = 4'b0111; // x=86, y=43
        pixel_data[43][87] = 4'b0111; // x=87, y=43
        pixel_data[43][88] = 4'b0000; // x=88, y=43
        pixel_data[43][89] = 4'b0000; // x=89, y=43
        pixel_data[43][90] = 4'b0000; // x=90, y=43
        pixel_data[43][91] = 4'b0000; // x=91, y=43
        pixel_data[43][92] = 4'b0000; // x=92, y=43
        pixel_data[43][93] = 4'b0111; // x=93, y=43
        pixel_data[43][94] = 4'b0111; // x=94, y=43
        pixel_data[43][95] = 4'b0111; // x=95, y=43
        pixel_data[43][96] = 4'b0111; // x=96, y=43
        pixel_data[43][97] = 4'b0111; // x=97, y=43
        pixel_data[43][98] = 4'b0111; // x=98, y=43
        pixel_data[43][99] = 4'b0111; // x=99, y=43
        pixel_data[43][100] = 4'b0111; // x=100, y=43
        pixel_data[43][101] = 4'b0111; // x=101, y=43
        pixel_data[43][102] = 4'b0111; // x=102, y=43
        pixel_data[43][103] = 4'b0111; // x=103, y=43
        pixel_data[43][104] = 4'b0111; // x=104, y=43
        pixel_data[43][105] = 4'b0111; // x=105, y=43
        pixel_data[43][106] = 4'b0111; // x=106, y=43
        pixel_data[43][107] = 4'b0111; // x=107, y=43
        pixel_data[43][108] = 4'b0111; // x=108, y=43
        pixel_data[43][109] = 4'b0111; // x=109, y=43
        pixel_data[43][110] = 4'b0111; // x=110, y=43
        pixel_data[43][111] = 4'b0111; // x=111, y=43
        pixel_data[43][112] = 4'b0000; // x=112, y=43
        pixel_data[43][113] = 4'b0000; // x=113, y=43
        pixel_data[43][114] = 4'b0111; // x=114, y=43
        pixel_data[43][115] = 4'b0111; // x=115, y=43
        pixel_data[43][116] = 4'b0111; // x=116, y=43
        pixel_data[43][117] = 4'b0111; // x=117, y=43
        pixel_data[43][118] = 4'b0000; // x=118, y=43
        pixel_data[43][119] = 4'b0000; // x=119, y=43
        pixel_data[43][120] = 4'b0111; // x=120, y=43
        pixel_data[43][121] = 4'b0111; // x=121, y=43
        pixel_data[43][122] = 4'b0111; // x=122, y=43
        pixel_data[43][123] = 4'b0111; // x=123, y=43
        pixel_data[43][124] = 4'b0111; // x=124, y=43
        pixel_data[43][125] = 4'b0111; // x=125, y=43
        pixel_data[43][126] = 4'b0111; // x=126, y=43
        pixel_data[43][127] = 4'b0111; // x=127, y=43
        pixel_data[43][128] = 4'b0111; // x=128, y=43
        pixel_data[43][129] = 4'b0111; // x=129, y=43
        pixel_data[43][130] = 4'b0111; // x=130, y=43
        pixel_data[43][131] = 4'b0111; // x=131, y=43
        pixel_data[43][132] = 4'b0111; // x=132, y=43
        pixel_data[43][133] = 4'b0111; // x=133, y=43
        pixel_data[43][134] = 4'b0111; // x=134, y=43
        pixel_data[43][135] = 4'b0111; // x=135, y=43
        pixel_data[43][136] = 4'b0111; // x=136, y=43
        pixel_data[43][137] = 4'b0111; // x=137, y=43
        pixel_data[43][138] = 4'b0111; // x=138, y=43
        pixel_data[43][139] = 4'b0111; // x=139, y=43
        pixel_data[43][140] = 4'b0111; // x=140, y=43
        pixel_data[43][141] = 4'b0111; // x=141, y=43
        pixel_data[43][142] = 4'b0111; // x=142, y=43
        pixel_data[43][143] = 4'b0111; // x=143, y=43
        pixel_data[43][144] = 4'b0111; // x=144, y=43
        pixel_data[43][145] = 4'b0111; // x=145, y=43
        pixel_data[43][146] = 4'b0111; // x=146, y=43
        pixel_data[43][147] = 4'b0000; // x=147, y=43
        pixel_data[43][148] = 4'b0111; // x=148, y=43
        pixel_data[43][149] = 4'b0111; // x=149, y=43
        pixel_data[43][150] = 4'b0111; // x=150, y=43
        pixel_data[43][151] = 4'b0111; // x=151, y=43
        pixel_data[43][152] = 4'b0111; // x=152, y=43
        pixel_data[43][153] = 4'b0111; // x=153, y=43
        pixel_data[43][154] = 4'b0111; // x=154, y=43
        pixel_data[43][155] = 4'b0111; // x=155, y=43
        pixel_data[43][156] = 4'b0111; // x=156, y=43
        pixel_data[43][157] = 4'b0111; // x=157, y=43
        pixel_data[43][158] = 4'b0111; // x=158, y=43
        pixel_data[43][159] = 4'b0111; // x=159, y=43
        pixel_data[43][160] = 4'b0111; // x=160, y=43
        pixel_data[43][161] = 4'b0111; // x=161, y=43
        pixel_data[43][162] = 4'b0111; // x=162, y=43
        pixel_data[43][163] = 4'b0111; // x=163, y=43
        pixel_data[43][164] = 4'b0111; // x=164, y=43
        pixel_data[43][165] = 4'b0111; // x=165, y=43
        pixel_data[43][166] = 4'b0111; // x=166, y=43
        pixel_data[43][167] = 4'b0111; // x=167, y=43
        pixel_data[43][168] = 4'b0111; // x=168, y=43
        pixel_data[43][169] = 4'b0111; // x=169, y=43
        pixel_data[43][170] = 4'b0111; // x=170, y=43
        pixel_data[43][171] = 4'b0111; // x=171, y=43
        pixel_data[43][172] = 4'b0111; // x=172, y=43
        pixel_data[43][173] = 4'b0111; // x=173, y=43
        pixel_data[43][174] = 4'b0111; // x=174, y=43
        pixel_data[43][175] = 4'b0111; // x=175, y=43
        pixel_data[43][176] = 4'b0111; // x=176, y=43
        pixel_data[43][177] = 4'b0111; // x=177, y=43
        pixel_data[43][178] = 4'b0111; // x=178, y=43
        pixel_data[43][179] = 4'b0111; // x=179, y=43
        pixel_data[44][0] = 4'b0111; // x=0, y=44
        pixel_data[44][1] = 4'b0111; // x=1, y=44
        pixel_data[44][2] = 4'b0111; // x=2, y=44
        pixel_data[44][3] = 4'b0111; // x=3, y=44
        pixel_data[44][4] = 4'b0111; // x=4, y=44
        pixel_data[44][5] = 4'b0111; // x=5, y=44
        pixel_data[44][6] = 4'b0111; // x=6, y=44
        pixel_data[44][7] = 4'b0111; // x=7, y=44
        pixel_data[44][8] = 4'b0111; // x=8, y=44
        pixel_data[44][9] = 4'b0111; // x=9, y=44
        pixel_data[44][10] = 4'b0111; // x=10, y=44
        pixel_data[44][11] = 4'b0111; // x=11, y=44
        pixel_data[44][12] = 4'b0111; // x=12, y=44
        pixel_data[44][13] = 4'b0111; // x=13, y=44
        pixel_data[44][14] = 4'b0111; // x=14, y=44
        pixel_data[44][15] = 4'b0111; // x=15, y=44
        pixel_data[44][16] = 4'b0111; // x=16, y=44
        pixel_data[44][17] = 4'b0111; // x=17, y=44
        pixel_data[44][18] = 4'b0111; // x=18, y=44
        pixel_data[44][19] = 4'b0111; // x=19, y=44
        pixel_data[44][20] = 4'b0111; // x=20, y=44
        pixel_data[44][21] = 4'b0111; // x=21, y=44
        pixel_data[44][22] = 4'b0111; // x=22, y=44
        pixel_data[44][23] = 4'b0111; // x=23, y=44
        pixel_data[44][24] = 4'b0111; // x=24, y=44
        pixel_data[44][25] = 4'b0111; // x=25, y=44
        pixel_data[44][26] = 4'b0111; // x=26, y=44
        pixel_data[44][27] = 4'b0111; // x=27, y=44
        pixel_data[44][28] = 4'b0111; // x=28, y=44
        pixel_data[44][29] = 4'b0111; // x=29, y=44
        pixel_data[44][30] = 4'b0111; // x=30, y=44
        pixel_data[44][31] = 4'b0111; // x=31, y=44
        pixel_data[44][32] = 4'b0111; // x=32, y=44
        pixel_data[44][33] = 4'b0111; // x=33, y=44
        pixel_data[44][34] = 4'b0111; // x=34, y=44
        pixel_data[44][35] = 4'b0111; // x=35, y=44
        pixel_data[44][36] = 4'b0111; // x=36, y=44
        pixel_data[44][37] = 4'b0111; // x=37, y=44
        pixel_data[44][38] = 4'b0111; // x=38, y=44
        pixel_data[44][39] = 4'b0111; // x=39, y=44
        pixel_data[44][40] = 4'b0111; // x=40, y=44
        pixel_data[44][41] = 4'b0111; // x=41, y=44
        pixel_data[44][42] = 4'b0111; // x=42, y=44
        pixel_data[44][43] = 4'b0111; // x=43, y=44
        pixel_data[44][44] = 4'b0111; // x=44, y=44
        pixel_data[44][45] = 4'b0111; // x=45, y=44
        pixel_data[44][46] = 4'b0111; // x=46, y=44
        pixel_data[44][47] = 4'b0111; // x=47, y=44
        pixel_data[44][48] = 4'b0111; // x=48, y=44
        pixel_data[44][49] = 4'b0111; // x=49, y=44
        pixel_data[44][50] = 4'b0111; // x=50, y=44
        pixel_data[44][51] = 4'b0111; // x=51, y=44
        pixel_data[44][52] = 4'b0111; // x=52, y=44
        pixel_data[44][53] = 4'b0111; // x=53, y=44
        pixel_data[44][54] = 4'b0111; // x=54, y=44
        pixel_data[44][55] = 4'b0111; // x=55, y=44
        pixel_data[44][56] = 4'b0111; // x=56, y=44
        pixel_data[44][57] = 4'b0111; // x=57, y=44
        pixel_data[44][58] = 4'b0111; // x=58, y=44
        pixel_data[44][59] = 4'b0111; // x=59, y=44
        pixel_data[44][60] = 4'b0111; // x=60, y=44
        pixel_data[44][61] = 4'b0111; // x=61, y=44
        pixel_data[44][62] = 4'b0111; // x=62, y=44
        pixel_data[44][63] = 4'b0111; // x=63, y=44
        pixel_data[44][64] = 4'b0111; // x=64, y=44
        pixel_data[44][65] = 4'b0111; // x=65, y=44
        pixel_data[44][66] = 4'b0111; // x=66, y=44
        pixel_data[44][67] = 4'b0111; // x=67, y=44
        pixel_data[44][68] = 4'b0111; // x=68, y=44
        pixel_data[44][69] = 4'b0111; // x=69, y=44
        pixel_data[44][70] = 4'b0111; // x=70, y=44
        pixel_data[44][71] = 4'b0111; // x=71, y=44
        pixel_data[44][72] = 4'b0111; // x=72, y=44
        pixel_data[44][73] = 4'b0111; // x=73, y=44
        pixel_data[44][74] = 4'b0111; // x=74, y=44
        pixel_data[44][75] = 4'b0111; // x=75, y=44
        pixel_data[44][76] = 4'b0111; // x=76, y=44
        pixel_data[44][77] = 4'b0111; // x=77, y=44
        pixel_data[44][78] = 4'b0111; // x=78, y=44
        pixel_data[44][79] = 4'b0111; // x=79, y=44
        pixel_data[44][80] = 4'b0111; // x=80, y=44
        pixel_data[44][81] = 4'b0111; // x=81, y=44
        pixel_data[44][82] = 4'b0111; // x=82, y=44
        pixel_data[44][83] = 4'b0111; // x=83, y=44
        pixel_data[44][84] = 4'b0111; // x=84, y=44
        pixel_data[44][85] = 4'b0111; // x=85, y=44
        pixel_data[44][86] = 4'b0111; // x=86, y=44
        pixel_data[44][87] = 4'b0111; // x=87, y=44
        pixel_data[44][88] = 4'b0111; // x=88, y=44
        pixel_data[44][89] = 4'b0111; // x=89, y=44
        pixel_data[44][90] = 4'b0111; // x=90, y=44
        pixel_data[44][91] = 4'b0111; // x=91, y=44
        pixel_data[44][92] = 4'b0111; // x=92, y=44
        pixel_data[44][93] = 4'b0111; // x=93, y=44
        pixel_data[44][94] = 4'b0111; // x=94, y=44
        pixel_data[44][95] = 4'b0111; // x=95, y=44
        pixel_data[44][96] = 4'b0111; // x=96, y=44
        pixel_data[44][97] = 4'b0111; // x=97, y=44
        pixel_data[44][98] = 4'b0111; // x=98, y=44
        pixel_data[44][99] = 4'b0111; // x=99, y=44
        pixel_data[44][100] = 4'b0111; // x=100, y=44
        pixel_data[44][101] = 4'b0111; // x=101, y=44
        pixel_data[44][102] = 4'b0111; // x=102, y=44
        pixel_data[44][103] = 4'b0111; // x=103, y=44
        pixel_data[44][104] = 4'b0111; // x=104, y=44
        pixel_data[44][105] = 4'b0111; // x=105, y=44
        pixel_data[44][106] = 4'b0111; // x=106, y=44
        pixel_data[44][107] = 4'b0111; // x=107, y=44
        pixel_data[44][108] = 4'b0111; // x=108, y=44
        pixel_data[44][109] = 4'b0111; // x=109, y=44
        pixel_data[44][110] = 4'b0111; // x=110, y=44
        pixel_data[44][111] = 4'b0111; // x=111, y=44
        pixel_data[44][112] = 4'b0111; // x=112, y=44
        pixel_data[44][113] = 4'b0111; // x=113, y=44
        pixel_data[44][114] = 4'b0111; // x=114, y=44
        pixel_data[44][115] = 4'b0111; // x=115, y=44
        pixel_data[44][116] = 4'b0111; // x=116, y=44
        pixel_data[44][117] = 4'b0111; // x=117, y=44
        pixel_data[44][118] = 4'b0111; // x=118, y=44
        pixel_data[44][119] = 4'b0111; // x=119, y=44
        pixel_data[44][120] = 4'b0111; // x=120, y=44
        pixel_data[44][121] = 4'b0111; // x=121, y=44
        pixel_data[44][122] = 4'b0111; // x=122, y=44
        pixel_data[44][123] = 4'b0111; // x=123, y=44
        pixel_data[44][124] = 4'b0111; // x=124, y=44
        pixel_data[44][125] = 4'b0111; // x=125, y=44
        pixel_data[44][126] = 4'b0111; // x=126, y=44
        pixel_data[44][127] = 4'b0111; // x=127, y=44
        pixel_data[44][128] = 4'b0111; // x=128, y=44
        pixel_data[44][129] = 4'b0111; // x=129, y=44
        pixel_data[44][130] = 4'b0111; // x=130, y=44
        pixel_data[44][131] = 4'b0111; // x=131, y=44
        pixel_data[44][132] = 4'b0111; // x=132, y=44
        pixel_data[44][133] = 4'b0111; // x=133, y=44
        pixel_data[44][134] = 4'b0111; // x=134, y=44
        pixel_data[44][135] = 4'b0111; // x=135, y=44
        pixel_data[44][136] = 4'b0111; // x=136, y=44
        pixel_data[44][137] = 4'b0111; // x=137, y=44
        pixel_data[44][138] = 4'b0111; // x=138, y=44
        pixel_data[44][139] = 4'b0111; // x=139, y=44
        pixel_data[44][140] = 4'b0111; // x=140, y=44
        pixel_data[44][141] = 4'b0111; // x=141, y=44
        pixel_data[44][142] = 4'b0111; // x=142, y=44
        pixel_data[44][143] = 4'b0111; // x=143, y=44
        pixel_data[44][144] = 4'b0111; // x=144, y=44
        pixel_data[44][145] = 4'b0111; // x=145, y=44
        pixel_data[44][146] = 4'b0111; // x=146, y=44
        pixel_data[44][147] = 4'b0111; // x=147, y=44
        pixel_data[44][148] = 4'b0111; // x=148, y=44
        pixel_data[44][149] = 4'b0111; // x=149, y=44
        pixel_data[44][150] = 4'b0111; // x=150, y=44
        pixel_data[44][151] = 4'b0111; // x=151, y=44
        pixel_data[44][152] = 4'b0111; // x=152, y=44
        pixel_data[44][153] = 4'b0111; // x=153, y=44
        pixel_data[44][154] = 4'b0111; // x=154, y=44
        pixel_data[44][155] = 4'b0111; // x=155, y=44
        pixel_data[44][156] = 4'b0111; // x=156, y=44
        pixel_data[44][157] = 4'b0111; // x=157, y=44
        pixel_data[44][158] = 4'b0111; // x=158, y=44
        pixel_data[44][159] = 4'b0111; // x=159, y=44
        pixel_data[44][160] = 4'b0111; // x=160, y=44
        pixel_data[44][161] = 4'b0111; // x=161, y=44
        pixel_data[44][162] = 4'b0111; // x=162, y=44
        pixel_data[44][163] = 4'b0111; // x=163, y=44
        pixel_data[44][164] = 4'b0111; // x=164, y=44
        pixel_data[44][165] = 4'b0111; // x=165, y=44
        pixel_data[44][166] = 4'b0111; // x=166, y=44
        pixel_data[44][167] = 4'b0111; // x=167, y=44
        pixel_data[44][168] = 4'b0111; // x=168, y=44
        pixel_data[44][169] = 4'b0111; // x=169, y=44
        pixel_data[44][170] = 4'b0111; // x=170, y=44
        pixel_data[44][171] = 4'b0111; // x=171, y=44
        pixel_data[44][172] = 4'b0111; // x=172, y=44
        pixel_data[44][173] = 4'b0111; // x=173, y=44
        pixel_data[44][174] = 4'b0111; // x=174, y=44
        pixel_data[44][175] = 4'b0111; // x=175, y=44
        pixel_data[44][176] = 4'b0111; // x=176, y=44
        pixel_data[44][177] = 4'b0111; // x=177, y=44
        pixel_data[44][178] = 4'b0111; // x=178, y=44
        pixel_data[44][179] = 4'b0111; // x=179, y=44
        pixel_data[45][0] = 4'b0111; // x=0, y=45
        pixel_data[45][1] = 4'b0111; // x=1, y=45
        pixel_data[45][2] = 4'b0111; // x=2, y=45
        pixel_data[45][3] = 4'b0111; // x=3, y=45
        pixel_data[45][4] = 4'b0111; // x=4, y=45
        pixel_data[45][5] = 4'b0111; // x=5, y=45
        pixel_data[45][6] = 4'b0111; // x=6, y=45
        pixel_data[45][7] = 4'b0111; // x=7, y=45
        pixel_data[45][8] = 4'b0111; // x=8, y=45
        pixel_data[45][9] = 4'b0111; // x=9, y=45
        pixel_data[45][10] = 4'b0111; // x=10, y=45
        pixel_data[45][11] = 4'b0111; // x=11, y=45
        pixel_data[45][12] = 4'b0111; // x=12, y=45
        pixel_data[45][13] = 4'b0111; // x=13, y=45
        pixel_data[45][14] = 4'b0111; // x=14, y=45
        pixel_data[45][15] = 4'b0111; // x=15, y=45
        pixel_data[45][16] = 4'b0111; // x=16, y=45
        pixel_data[45][17] = 4'b0111; // x=17, y=45
        pixel_data[45][18] = 4'b0111; // x=18, y=45
        pixel_data[45][19] = 4'b0111; // x=19, y=45
        pixel_data[45][20] = 4'b0111; // x=20, y=45
        pixel_data[45][21] = 4'b0111; // x=21, y=45
        pixel_data[45][22] = 4'b0111; // x=22, y=45
        pixel_data[45][23] = 4'b0111; // x=23, y=45
        pixel_data[45][24] = 4'b0111; // x=24, y=45
        pixel_data[45][25] = 4'b0111; // x=25, y=45
        pixel_data[45][26] = 4'b0111; // x=26, y=45
        pixel_data[45][27] = 4'b0111; // x=27, y=45
        pixel_data[45][28] = 4'b0111; // x=28, y=45
        pixel_data[45][29] = 4'b0111; // x=29, y=45
        pixel_data[45][30] = 4'b0111; // x=30, y=45
        pixel_data[45][31] = 4'b0111; // x=31, y=45
        pixel_data[45][32] = 4'b0111; // x=32, y=45
        pixel_data[45][33] = 4'b0111; // x=33, y=45
        pixel_data[45][34] = 4'b0111; // x=34, y=45
        pixel_data[45][35] = 4'b0111; // x=35, y=45
        pixel_data[45][36] = 4'b0111; // x=36, y=45
        pixel_data[45][37] = 4'b0111; // x=37, y=45
        pixel_data[45][38] = 4'b0111; // x=38, y=45
        pixel_data[45][39] = 4'b0111; // x=39, y=45
        pixel_data[45][40] = 4'b0111; // x=40, y=45
        pixel_data[45][41] = 4'b0111; // x=41, y=45
        pixel_data[45][42] = 4'b0111; // x=42, y=45
        pixel_data[45][43] = 4'b0111; // x=43, y=45
        pixel_data[45][44] = 4'b0111; // x=44, y=45
        pixel_data[45][45] = 4'b0111; // x=45, y=45
        pixel_data[45][46] = 4'b0111; // x=46, y=45
        pixel_data[45][47] = 4'b0111; // x=47, y=45
        pixel_data[45][48] = 4'b0111; // x=48, y=45
        pixel_data[45][49] = 4'b0111; // x=49, y=45
        pixel_data[45][50] = 4'b0111; // x=50, y=45
        pixel_data[45][51] = 4'b0111; // x=51, y=45
        pixel_data[45][52] = 4'b0111; // x=52, y=45
        pixel_data[45][53] = 4'b0111; // x=53, y=45
        pixel_data[45][54] = 4'b0111; // x=54, y=45
        pixel_data[45][55] = 4'b0111; // x=55, y=45
        pixel_data[45][56] = 4'b0111; // x=56, y=45
        pixel_data[45][57] = 4'b0111; // x=57, y=45
        pixel_data[45][58] = 4'b0111; // x=58, y=45
        pixel_data[45][59] = 4'b0111; // x=59, y=45
        pixel_data[45][60] = 4'b0111; // x=60, y=45
        pixel_data[45][61] = 4'b0111; // x=61, y=45
        pixel_data[45][62] = 4'b0111; // x=62, y=45
        pixel_data[45][63] = 4'b0111; // x=63, y=45
        pixel_data[45][64] = 4'b0111; // x=64, y=45
        pixel_data[45][65] = 4'b0111; // x=65, y=45
        pixel_data[45][66] = 4'b0111; // x=66, y=45
        pixel_data[45][67] = 4'b0111; // x=67, y=45
        pixel_data[45][68] = 4'b0111; // x=68, y=45
        pixel_data[45][69] = 4'b0111; // x=69, y=45
        pixel_data[45][70] = 4'b0111; // x=70, y=45
        pixel_data[45][71] = 4'b0111; // x=71, y=45
        pixel_data[45][72] = 4'b0111; // x=72, y=45
        pixel_data[45][73] = 4'b0111; // x=73, y=45
        pixel_data[45][74] = 4'b0111; // x=74, y=45
        pixel_data[45][75] = 4'b0111; // x=75, y=45
        pixel_data[45][76] = 4'b0111; // x=76, y=45
        pixel_data[45][77] = 4'b0111; // x=77, y=45
        pixel_data[45][78] = 4'b0111; // x=78, y=45
        pixel_data[45][79] = 4'b0111; // x=79, y=45
        pixel_data[45][80] = 4'b0111; // x=80, y=45
        pixel_data[45][81] = 4'b0111; // x=81, y=45
        pixel_data[45][82] = 4'b0111; // x=82, y=45
        pixel_data[45][83] = 4'b0111; // x=83, y=45
        pixel_data[45][84] = 4'b0111; // x=84, y=45
        pixel_data[45][85] = 4'b0111; // x=85, y=45
        pixel_data[45][86] = 4'b0111; // x=86, y=45
        pixel_data[45][87] = 4'b0111; // x=87, y=45
        pixel_data[45][88] = 4'b0111; // x=88, y=45
        pixel_data[45][89] = 4'b0111; // x=89, y=45
        pixel_data[45][90] = 4'b0111; // x=90, y=45
        pixel_data[45][91] = 4'b0111; // x=91, y=45
        pixel_data[45][92] = 4'b0111; // x=92, y=45
        pixel_data[45][93] = 4'b0111; // x=93, y=45
        pixel_data[45][94] = 4'b0111; // x=94, y=45
        pixel_data[45][95] = 4'b0111; // x=95, y=45
        pixel_data[45][96] = 4'b0111; // x=96, y=45
        pixel_data[45][97] = 4'b0111; // x=97, y=45
        pixel_data[45][98] = 4'b0111; // x=98, y=45
        pixel_data[45][99] = 4'b0111; // x=99, y=45
        pixel_data[45][100] = 4'b0111; // x=100, y=45
        pixel_data[45][101] = 4'b0111; // x=101, y=45
        pixel_data[45][102] = 4'b0111; // x=102, y=45
        pixel_data[45][103] = 4'b0111; // x=103, y=45
        pixel_data[45][104] = 4'b0111; // x=104, y=45
        pixel_data[45][105] = 4'b0111; // x=105, y=45
        pixel_data[45][106] = 4'b0111; // x=106, y=45
        pixel_data[45][107] = 4'b0111; // x=107, y=45
        pixel_data[45][108] = 4'b0111; // x=108, y=45
        pixel_data[45][109] = 4'b0111; // x=109, y=45
        pixel_data[45][110] = 4'b0111; // x=110, y=45
        pixel_data[45][111] = 4'b0111; // x=111, y=45
        pixel_data[45][112] = 4'b0111; // x=112, y=45
        pixel_data[45][113] = 4'b0111; // x=113, y=45
        pixel_data[45][114] = 4'b0111; // x=114, y=45
        pixel_data[45][115] = 4'b0111; // x=115, y=45
        pixel_data[45][116] = 4'b0111; // x=116, y=45
        pixel_data[45][117] = 4'b0111; // x=117, y=45
        pixel_data[45][118] = 4'b0111; // x=118, y=45
        pixel_data[45][119] = 4'b0111; // x=119, y=45
        pixel_data[45][120] = 4'b0111; // x=120, y=45
        pixel_data[45][121] = 4'b0111; // x=121, y=45
        pixel_data[45][122] = 4'b0111; // x=122, y=45
        pixel_data[45][123] = 4'b0111; // x=123, y=45
        pixel_data[45][124] = 4'b0111; // x=124, y=45
        pixel_data[45][125] = 4'b0111; // x=125, y=45
        pixel_data[45][126] = 4'b0111; // x=126, y=45
        pixel_data[45][127] = 4'b0111; // x=127, y=45
        pixel_data[45][128] = 4'b0111; // x=128, y=45
        pixel_data[45][129] = 4'b0111; // x=129, y=45
        pixel_data[45][130] = 4'b0111; // x=130, y=45
        pixel_data[45][131] = 4'b0111; // x=131, y=45
        pixel_data[45][132] = 4'b0111; // x=132, y=45
        pixel_data[45][133] = 4'b0111; // x=133, y=45
        pixel_data[45][134] = 4'b0111; // x=134, y=45
        pixel_data[45][135] = 4'b0111; // x=135, y=45
        pixel_data[45][136] = 4'b0111; // x=136, y=45
        pixel_data[45][137] = 4'b0111; // x=137, y=45
        pixel_data[45][138] = 4'b0111; // x=138, y=45
        pixel_data[45][139] = 4'b0111; // x=139, y=45
        pixel_data[45][140] = 4'b0111; // x=140, y=45
        pixel_data[45][141] = 4'b0111; // x=141, y=45
        pixel_data[45][142] = 4'b0111; // x=142, y=45
        pixel_data[45][143] = 4'b0111; // x=143, y=45
        pixel_data[45][144] = 4'b0111; // x=144, y=45
        pixel_data[45][145] = 4'b0111; // x=145, y=45
        pixel_data[45][146] = 4'b0111; // x=146, y=45
        pixel_data[45][147] = 4'b0111; // x=147, y=45
        pixel_data[45][148] = 4'b0111; // x=148, y=45
        pixel_data[45][149] = 4'b0111; // x=149, y=45
        pixel_data[45][150] = 4'b0111; // x=150, y=45
        pixel_data[45][151] = 4'b0111; // x=151, y=45
        pixel_data[45][152] = 4'b0111; // x=152, y=45
        pixel_data[45][153] = 4'b0111; // x=153, y=45
        pixel_data[45][154] = 4'b0111; // x=154, y=45
        pixel_data[45][155] = 4'b0111; // x=155, y=45
        pixel_data[45][156] = 4'b0111; // x=156, y=45
        pixel_data[45][157] = 4'b0111; // x=157, y=45
        pixel_data[45][158] = 4'b0111; // x=158, y=45
        pixel_data[45][159] = 4'b0111; // x=159, y=45
        pixel_data[45][160] = 4'b0111; // x=160, y=45
        pixel_data[45][161] = 4'b0111; // x=161, y=45
        pixel_data[45][162] = 4'b0111; // x=162, y=45
        pixel_data[45][163] = 4'b0111; // x=163, y=45
        pixel_data[45][164] = 4'b0111; // x=164, y=45
        pixel_data[45][165] = 4'b0111; // x=165, y=45
        pixel_data[45][166] = 4'b0111; // x=166, y=45
        pixel_data[45][167] = 4'b0111; // x=167, y=45
        pixel_data[45][168] = 4'b0111; // x=168, y=45
        pixel_data[45][169] = 4'b0111; // x=169, y=45
        pixel_data[45][170] = 4'b0111; // x=170, y=45
        pixel_data[45][171] = 4'b0111; // x=171, y=45
        pixel_data[45][172] = 4'b0111; // x=172, y=45
        pixel_data[45][173] = 4'b0111; // x=173, y=45
        pixel_data[45][174] = 4'b0111; // x=174, y=45
        pixel_data[45][175] = 4'b0111; // x=175, y=45
        pixel_data[45][176] = 4'b0111; // x=176, y=45
        pixel_data[45][177] = 4'b0111; // x=177, y=45
        pixel_data[45][178] = 4'b0111; // x=178, y=45
        pixel_data[45][179] = 4'b0111; // x=179, y=45
        pixel_data[46][0] = 4'b0111; // x=0, y=46
        pixel_data[46][1] = 4'b0111; // x=1, y=46
        pixel_data[46][2] = 4'b0111; // x=2, y=46
        pixel_data[46][3] = 4'b0111; // x=3, y=46
        pixel_data[46][4] = 4'b0111; // x=4, y=46
        pixel_data[46][5] = 4'b0111; // x=5, y=46
        pixel_data[46][6] = 4'b0111; // x=6, y=46
        pixel_data[46][7] = 4'b0111; // x=7, y=46
        pixel_data[46][8] = 4'b0111; // x=8, y=46
        pixel_data[46][9] = 4'b0111; // x=9, y=46
        pixel_data[46][10] = 4'b0111; // x=10, y=46
        pixel_data[46][11] = 4'b0111; // x=11, y=46
        pixel_data[46][12] = 4'b0111; // x=12, y=46
        pixel_data[46][13] = 4'b0111; // x=13, y=46
        pixel_data[46][14] = 4'b0111; // x=14, y=46
        pixel_data[46][15] = 4'b0111; // x=15, y=46
        pixel_data[46][16] = 4'b0111; // x=16, y=46
        pixel_data[46][17] = 4'b0111; // x=17, y=46
        pixel_data[46][18] = 4'b0111; // x=18, y=46
        pixel_data[46][19] = 4'b0111; // x=19, y=46
        pixel_data[46][20] = 4'b0111; // x=20, y=46
        pixel_data[46][21] = 4'b0111; // x=21, y=46
        pixel_data[46][22] = 4'b0111; // x=22, y=46
        pixel_data[46][23] = 4'b0111; // x=23, y=46
        pixel_data[46][24] = 4'b0111; // x=24, y=46
        pixel_data[46][25] = 4'b0111; // x=25, y=46
        pixel_data[46][26] = 4'b0111; // x=26, y=46
        pixel_data[46][27] = 4'b0111; // x=27, y=46
        pixel_data[46][28] = 4'b0111; // x=28, y=46
        pixel_data[46][29] = 4'b0111; // x=29, y=46
        pixel_data[46][30] = 4'b0111; // x=30, y=46
        pixel_data[46][31] = 4'b0111; // x=31, y=46
        pixel_data[46][32] = 4'b0111; // x=32, y=46
        pixel_data[46][33] = 4'b0111; // x=33, y=46
        pixel_data[46][34] = 4'b0111; // x=34, y=46
        pixel_data[46][35] = 4'b0111; // x=35, y=46
        pixel_data[46][36] = 4'b0111; // x=36, y=46
        pixel_data[46][37] = 4'b0111; // x=37, y=46
        pixel_data[46][38] = 4'b0111; // x=38, y=46
        pixel_data[46][39] = 4'b0111; // x=39, y=46
        pixel_data[46][40] = 4'b0111; // x=40, y=46
        pixel_data[46][41] = 4'b0111; // x=41, y=46
        pixel_data[46][42] = 4'b0111; // x=42, y=46
        pixel_data[46][43] = 4'b0111; // x=43, y=46
        pixel_data[46][44] = 4'b0111; // x=44, y=46
        pixel_data[46][45] = 4'b0111; // x=45, y=46
        pixel_data[46][46] = 4'b0111; // x=46, y=46
        pixel_data[46][47] = 4'b0111; // x=47, y=46
        pixel_data[46][48] = 4'b0111; // x=48, y=46
        pixel_data[46][49] = 4'b0111; // x=49, y=46
        pixel_data[46][50] = 4'b0111; // x=50, y=46
        pixel_data[46][51] = 4'b0111; // x=51, y=46
        pixel_data[46][52] = 4'b0111; // x=52, y=46
        pixel_data[46][53] = 4'b0111; // x=53, y=46
        pixel_data[46][54] = 4'b0111; // x=54, y=46
        pixel_data[46][55] = 4'b0111; // x=55, y=46
        pixel_data[46][56] = 4'b0111; // x=56, y=46
        pixel_data[46][57] = 4'b0111; // x=57, y=46
        pixel_data[46][58] = 4'b0111; // x=58, y=46
        pixel_data[46][59] = 4'b0111; // x=59, y=46
        pixel_data[46][60] = 4'b0111; // x=60, y=46
        pixel_data[46][61] = 4'b0111; // x=61, y=46
        pixel_data[46][62] = 4'b0111; // x=62, y=46
        pixel_data[46][63] = 4'b0111; // x=63, y=46
        pixel_data[46][64] = 4'b0111; // x=64, y=46
        pixel_data[46][65] = 4'b0111; // x=65, y=46
        pixel_data[46][66] = 4'b0111; // x=66, y=46
        pixel_data[46][67] = 4'b0111; // x=67, y=46
        pixel_data[46][68] = 4'b0111; // x=68, y=46
        pixel_data[46][69] = 4'b0111; // x=69, y=46
        pixel_data[46][70] = 4'b0111; // x=70, y=46
        pixel_data[46][71] = 4'b0111; // x=71, y=46
        pixel_data[46][72] = 4'b0111; // x=72, y=46
        pixel_data[46][73] = 4'b0111; // x=73, y=46
        pixel_data[46][74] = 4'b0111; // x=74, y=46
        pixel_data[46][75] = 4'b0111; // x=75, y=46
        pixel_data[46][76] = 4'b0111; // x=76, y=46
        pixel_data[46][77] = 4'b0111; // x=77, y=46
        pixel_data[46][78] = 4'b0111; // x=78, y=46
        pixel_data[46][79] = 4'b0111; // x=79, y=46
        pixel_data[46][80] = 4'b0111; // x=80, y=46
        pixel_data[46][81] = 4'b0111; // x=81, y=46
        pixel_data[46][82] = 4'b0111; // x=82, y=46
        pixel_data[46][83] = 4'b0111; // x=83, y=46
        pixel_data[46][84] = 4'b0111; // x=84, y=46
        pixel_data[46][85] = 4'b0111; // x=85, y=46
        pixel_data[46][86] = 4'b0111; // x=86, y=46
        pixel_data[46][87] = 4'b0111; // x=87, y=46
        pixel_data[46][88] = 4'b0111; // x=88, y=46
        pixel_data[46][89] = 4'b0111; // x=89, y=46
        pixel_data[46][90] = 4'b0111; // x=90, y=46
        pixel_data[46][91] = 4'b0111; // x=91, y=46
        pixel_data[46][92] = 4'b0111; // x=92, y=46
        pixel_data[46][93] = 4'b0111; // x=93, y=46
        pixel_data[46][94] = 4'b0111; // x=94, y=46
        pixel_data[46][95] = 4'b0111; // x=95, y=46
        pixel_data[46][96] = 4'b0111; // x=96, y=46
        pixel_data[46][97] = 4'b0111; // x=97, y=46
        pixel_data[46][98] = 4'b0111; // x=98, y=46
        pixel_data[46][99] = 4'b0111; // x=99, y=46
        pixel_data[46][100] = 4'b0111; // x=100, y=46
        pixel_data[46][101] = 4'b0111; // x=101, y=46
        pixel_data[46][102] = 4'b0111; // x=102, y=46
        pixel_data[46][103] = 4'b0111; // x=103, y=46
        pixel_data[46][104] = 4'b0111; // x=104, y=46
        pixel_data[46][105] = 4'b0111; // x=105, y=46
        pixel_data[46][106] = 4'b0111; // x=106, y=46
        pixel_data[46][107] = 4'b0111; // x=107, y=46
        pixel_data[46][108] = 4'b0111; // x=108, y=46
        pixel_data[46][109] = 4'b0111; // x=109, y=46
        pixel_data[46][110] = 4'b0111; // x=110, y=46
        pixel_data[46][111] = 4'b0111; // x=111, y=46
        pixel_data[46][112] = 4'b0111; // x=112, y=46
        pixel_data[46][113] = 4'b0111; // x=113, y=46
        pixel_data[46][114] = 4'b0111; // x=114, y=46
        pixel_data[46][115] = 4'b0111; // x=115, y=46
        pixel_data[46][116] = 4'b0111; // x=116, y=46
        pixel_data[46][117] = 4'b0111; // x=117, y=46
        pixel_data[46][118] = 4'b0111; // x=118, y=46
        pixel_data[46][119] = 4'b0111; // x=119, y=46
        pixel_data[46][120] = 4'b0111; // x=120, y=46
        pixel_data[46][121] = 4'b0111; // x=121, y=46
        pixel_data[46][122] = 4'b0111; // x=122, y=46
        pixel_data[46][123] = 4'b0111; // x=123, y=46
        pixel_data[46][124] = 4'b0111; // x=124, y=46
        pixel_data[46][125] = 4'b0111; // x=125, y=46
        pixel_data[46][126] = 4'b0111; // x=126, y=46
        pixel_data[46][127] = 4'b0111; // x=127, y=46
        pixel_data[46][128] = 4'b0111; // x=128, y=46
        pixel_data[46][129] = 4'b0111; // x=129, y=46
        pixel_data[46][130] = 4'b0111; // x=130, y=46
        pixel_data[46][131] = 4'b0111; // x=131, y=46
        pixel_data[46][132] = 4'b0111; // x=132, y=46
        pixel_data[46][133] = 4'b0111; // x=133, y=46
        pixel_data[46][134] = 4'b0111; // x=134, y=46
        pixel_data[46][135] = 4'b0111; // x=135, y=46
        pixel_data[46][136] = 4'b0111; // x=136, y=46
        pixel_data[46][137] = 4'b0111; // x=137, y=46
        pixel_data[46][138] = 4'b0111; // x=138, y=46
        pixel_data[46][139] = 4'b0111; // x=139, y=46
        pixel_data[46][140] = 4'b0111; // x=140, y=46
        pixel_data[46][141] = 4'b0111; // x=141, y=46
        pixel_data[46][142] = 4'b0111; // x=142, y=46
        pixel_data[46][143] = 4'b0111; // x=143, y=46
        pixel_data[46][144] = 4'b0111; // x=144, y=46
        pixel_data[46][145] = 4'b0111; // x=145, y=46
        pixel_data[46][146] = 4'b0111; // x=146, y=46
        pixel_data[46][147] = 4'b0111; // x=147, y=46
        pixel_data[46][148] = 4'b0111; // x=148, y=46
        pixel_data[46][149] = 4'b0111; // x=149, y=46
        pixel_data[46][150] = 4'b0111; // x=150, y=46
        pixel_data[46][151] = 4'b0111; // x=151, y=46
        pixel_data[46][152] = 4'b0111; // x=152, y=46
        pixel_data[46][153] = 4'b0111; // x=153, y=46
        pixel_data[46][154] = 4'b0111; // x=154, y=46
        pixel_data[46][155] = 4'b0111; // x=155, y=46
        pixel_data[46][156] = 4'b0111; // x=156, y=46
        pixel_data[46][157] = 4'b0111; // x=157, y=46
        pixel_data[46][158] = 4'b0111; // x=158, y=46
        pixel_data[46][159] = 4'b0111; // x=159, y=46
        pixel_data[46][160] = 4'b0111; // x=160, y=46
        pixel_data[46][161] = 4'b0111; // x=161, y=46
        pixel_data[46][162] = 4'b0111; // x=162, y=46
        pixel_data[46][163] = 4'b0111; // x=163, y=46
        pixel_data[46][164] = 4'b0111; // x=164, y=46
        pixel_data[46][165] = 4'b0111; // x=165, y=46
        pixel_data[46][166] = 4'b0111; // x=166, y=46
        pixel_data[46][167] = 4'b0111; // x=167, y=46
        pixel_data[46][168] = 4'b0111; // x=168, y=46
        pixel_data[46][169] = 4'b0111; // x=169, y=46
        pixel_data[46][170] = 4'b0111; // x=170, y=46
        pixel_data[46][171] = 4'b0111; // x=171, y=46
        pixel_data[46][172] = 4'b0111; // x=172, y=46
        pixel_data[46][173] = 4'b0111; // x=173, y=46
        pixel_data[46][174] = 4'b0111; // x=174, y=46
        pixel_data[46][175] = 4'b0111; // x=175, y=46
        pixel_data[46][176] = 4'b0111; // x=176, y=46
        pixel_data[46][177] = 4'b0111; // x=177, y=46
        pixel_data[46][178] = 4'b0111; // x=178, y=46
        pixel_data[46][179] = 4'b0111; // x=179, y=46
        pixel_data[47][0] = 4'b0111; // x=0, y=47
        pixel_data[47][1] = 4'b0111; // x=1, y=47
        pixel_data[47][2] = 4'b0111; // x=2, y=47
        pixel_data[47][3] = 4'b0111; // x=3, y=47
        pixel_data[47][4] = 4'b0111; // x=4, y=47
        pixel_data[47][5] = 4'b0111; // x=5, y=47
        pixel_data[47][6] = 4'b0111; // x=6, y=47
        pixel_data[47][7] = 4'b0111; // x=7, y=47
        pixel_data[47][8] = 4'b0111; // x=8, y=47
        pixel_data[47][9] = 4'b0111; // x=9, y=47
        pixel_data[47][10] = 4'b0111; // x=10, y=47
        pixel_data[47][11] = 4'b0111; // x=11, y=47
        pixel_data[47][12] = 4'b0111; // x=12, y=47
        pixel_data[47][13] = 4'b0111; // x=13, y=47
        pixel_data[47][14] = 4'b0111; // x=14, y=47
        pixel_data[47][15] = 4'b0111; // x=15, y=47
        pixel_data[47][16] = 4'b0111; // x=16, y=47
        pixel_data[47][17] = 4'b0111; // x=17, y=47
        pixel_data[47][18] = 4'b0111; // x=18, y=47
        pixel_data[47][19] = 4'b0111; // x=19, y=47
        pixel_data[47][20] = 4'b0111; // x=20, y=47
        pixel_data[47][21] = 4'b0111; // x=21, y=47
        pixel_data[47][22] = 4'b0111; // x=22, y=47
        pixel_data[47][23] = 4'b0111; // x=23, y=47
        pixel_data[47][24] = 4'b0111; // x=24, y=47
        pixel_data[47][25] = 4'b0111; // x=25, y=47
        pixel_data[47][26] = 4'b0111; // x=26, y=47
        pixel_data[47][27] = 4'b0111; // x=27, y=47
        pixel_data[47][28] = 4'b0111; // x=28, y=47
        pixel_data[47][29] = 4'b0111; // x=29, y=47
        pixel_data[47][30] = 4'b0111; // x=30, y=47
        pixel_data[47][31] = 4'b0111; // x=31, y=47
        pixel_data[47][32] = 4'b0111; // x=32, y=47
        pixel_data[47][33] = 4'b0111; // x=33, y=47
        pixel_data[47][34] = 4'b0111; // x=34, y=47
        pixel_data[47][35] = 4'b0111; // x=35, y=47
        pixel_data[47][36] = 4'b0111; // x=36, y=47
        pixel_data[47][37] = 4'b0111; // x=37, y=47
        pixel_data[47][38] = 4'b0111; // x=38, y=47
        pixel_data[47][39] = 4'b0111; // x=39, y=47
        pixel_data[47][40] = 4'b0111; // x=40, y=47
        pixel_data[47][41] = 4'b0111; // x=41, y=47
        pixel_data[47][42] = 4'b0111; // x=42, y=47
        pixel_data[47][43] = 4'b0111; // x=43, y=47
        pixel_data[47][44] = 4'b0111; // x=44, y=47
        pixel_data[47][45] = 4'b0111; // x=45, y=47
        pixel_data[47][46] = 4'b0111; // x=46, y=47
        pixel_data[47][47] = 4'b0111; // x=47, y=47
        pixel_data[47][48] = 4'b0111; // x=48, y=47
        pixel_data[47][49] = 4'b0111; // x=49, y=47
        pixel_data[47][50] = 4'b0111; // x=50, y=47
        pixel_data[47][51] = 4'b0111; // x=51, y=47
        pixel_data[47][52] = 4'b0111; // x=52, y=47
        pixel_data[47][53] = 4'b0111; // x=53, y=47
        pixel_data[47][54] = 4'b0111; // x=54, y=47
        pixel_data[47][55] = 4'b0111; // x=55, y=47
        pixel_data[47][56] = 4'b0111; // x=56, y=47
        pixel_data[47][57] = 4'b0111; // x=57, y=47
        pixel_data[47][58] = 4'b0111; // x=58, y=47
        pixel_data[47][59] = 4'b0111; // x=59, y=47
        pixel_data[47][60] = 4'b0111; // x=60, y=47
        pixel_data[47][61] = 4'b0111; // x=61, y=47
        pixel_data[47][62] = 4'b0111; // x=62, y=47
        pixel_data[47][63] = 4'b0111; // x=63, y=47
        pixel_data[47][64] = 4'b0111; // x=64, y=47
        pixel_data[47][65] = 4'b0111; // x=65, y=47
        pixel_data[47][66] = 4'b0111; // x=66, y=47
        pixel_data[47][67] = 4'b0111; // x=67, y=47
        pixel_data[47][68] = 4'b0111; // x=68, y=47
        pixel_data[47][69] = 4'b0111; // x=69, y=47
        pixel_data[47][70] = 4'b0111; // x=70, y=47
        pixel_data[47][71] = 4'b0111; // x=71, y=47
        pixel_data[47][72] = 4'b0111; // x=72, y=47
        pixel_data[47][73] = 4'b0111; // x=73, y=47
        pixel_data[47][74] = 4'b0111; // x=74, y=47
        pixel_data[47][75] = 4'b0111; // x=75, y=47
        pixel_data[47][76] = 4'b0111; // x=76, y=47
        pixel_data[47][77] = 4'b0111; // x=77, y=47
        pixel_data[47][78] = 4'b0111; // x=78, y=47
        pixel_data[47][79] = 4'b0111; // x=79, y=47
        pixel_data[47][80] = 4'b0111; // x=80, y=47
        pixel_data[47][81] = 4'b0111; // x=81, y=47
        pixel_data[47][82] = 4'b0111; // x=82, y=47
        pixel_data[47][83] = 4'b0111; // x=83, y=47
        pixel_data[47][84] = 4'b0111; // x=84, y=47
        pixel_data[47][85] = 4'b0111; // x=85, y=47
        pixel_data[47][86] = 4'b0111; // x=86, y=47
        pixel_data[47][87] = 4'b0111; // x=87, y=47
        pixel_data[47][88] = 4'b0111; // x=88, y=47
        pixel_data[47][89] = 4'b0111; // x=89, y=47
        pixel_data[47][90] = 4'b0111; // x=90, y=47
        pixel_data[47][91] = 4'b0111; // x=91, y=47
        pixel_data[47][92] = 4'b0111; // x=92, y=47
        pixel_data[47][93] = 4'b0111; // x=93, y=47
        pixel_data[47][94] = 4'b0111; // x=94, y=47
        pixel_data[47][95] = 4'b0111; // x=95, y=47
        pixel_data[47][96] = 4'b0111; // x=96, y=47
        pixel_data[47][97] = 4'b0111; // x=97, y=47
        pixel_data[47][98] = 4'b0111; // x=98, y=47
        pixel_data[47][99] = 4'b0111; // x=99, y=47
        pixel_data[47][100] = 4'b0111; // x=100, y=47
        pixel_data[47][101] = 4'b0111; // x=101, y=47
        pixel_data[47][102] = 4'b0111; // x=102, y=47
        pixel_data[47][103] = 4'b0111; // x=103, y=47
        pixel_data[47][104] = 4'b0111; // x=104, y=47
        pixel_data[47][105] = 4'b0111; // x=105, y=47
        pixel_data[47][106] = 4'b0111; // x=106, y=47
        pixel_data[47][107] = 4'b0111; // x=107, y=47
        pixel_data[47][108] = 4'b0111; // x=108, y=47
        pixel_data[47][109] = 4'b0111; // x=109, y=47
        pixel_data[47][110] = 4'b0111; // x=110, y=47
        pixel_data[47][111] = 4'b0111; // x=111, y=47
        pixel_data[47][112] = 4'b0111; // x=112, y=47
        pixel_data[47][113] = 4'b0111; // x=113, y=47
        pixel_data[47][114] = 4'b0111; // x=114, y=47
        pixel_data[47][115] = 4'b0111; // x=115, y=47
        pixel_data[47][116] = 4'b0111; // x=116, y=47
        pixel_data[47][117] = 4'b0111; // x=117, y=47
        pixel_data[47][118] = 4'b0111; // x=118, y=47
        pixel_data[47][119] = 4'b0111; // x=119, y=47
        pixel_data[47][120] = 4'b0111; // x=120, y=47
        pixel_data[47][121] = 4'b0111; // x=121, y=47
        pixel_data[47][122] = 4'b0111; // x=122, y=47
        pixel_data[47][123] = 4'b0111; // x=123, y=47
        pixel_data[47][124] = 4'b0111; // x=124, y=47
        pixel_data[47][125] = 4'b0111; // x=125, y=47
        pixel_data[47][126] = 4'b0111; // x=126, y=47
        pixel_data[47][127] = 4'b0111; // x=127, y=47
        pixel_data[47][128] = 4'b0111; // x=128, y=47
        pixel_data[47][129] = 4'b0111; // x=129, y=47
        pixel_data[47][130] = 4'b0111; // x=130, y=47
        pixel_data[47][131] = 4'b0111; // x=131, y=47
        pixel_data[47][132] = 4'b0111; // x=132, y=47
        pixel_data[47][133] = 4'b0111; // x=133, y=47
        pixel_data[47][134] = 4'b0111; // x=134, y=47
        pixel_data[47][135] = 4'b0111; // x=135, y=47
        pixel_data[47][136] = 4'b0111; // x=136, y=47
        pixel_data[47][137] = 4'b0111; // x=137, y=47
        pixel_data[47][138] = 4'b0111; // x=138, y=47
        pixel_data[47][139] = 4'b0111; // x=139, y=47
        pixel_data[47][140] = 4'b0111; // x=140, y=47
        pixel_data[47][141] = 4'b0111; // x=141, y=47
        pixel_data[47][142] = 4'b0111; // x=142, y=47
        pixel_data[47][143] = 4'b0111; // x=143, y=47
        pixel_data[47][144] = 4'b0111; // x=144, y=47
        pixel_data[47][145] = 4'b0111; // x=145, y=47
        pixel_data[47][146] = 4'b0111; // x=146, y=47
        pixel_data[47][147] = 4'b0111; // x=147, y=47
        pixel_data[47][148] = 4'b0111; // x=148, y=47
        pixel_data[47][149] = 4'b0111; // x=149, y=47
        pixel_data[47][150] = 4'b0111; // x=150, y=47
        pixel_data[47][151] = 4'b0111; // x=151, y=47
        pixel_data[47][152] = 4'b0111; // x=152, y=47
        pixel_data[47][153] = 4'b0111; // x=153, y=47
        pixel_data[47][154] = 4'b0111; // x=154, y=47
        pixel_data[47][155] = 4'b0111; // x=155, y=47
        pixel_data[47][156] = 4'b0111; // x=156, y=47
        pixel_data[47][157] = 4'b0111; // x=157, y=47
        pixel_data[47][158] = 4'b0111; // x=158, y=47
        pixel_data[47][159] = 4'b0111; // x=159, y=47
        pixel_data[47][160] = 4'b0111; // x=160, y=47
        pixel_data[47][161] = 4'b0111; // x=161, y=47
        pixel_data[47][162] = 4'b0111; // x=162, y=47
        pixel_data[47][163] = 4'b0111; // x=163, y=47
        pixel_data[47][164] = 4'b0111; // x=164, y=47
        pixel_data[47][165] = 4'b0111; // x=165, y=47
        pixel_data[47][166] = 4'b0111; // x=166, y=47
        pixel_data[47][167] = 4'b0111; // x=167, y=47
        pixel_data[47][168] = 4'b0111; // x=168, y=47
        pixel_data[47][169] = 4'b0111; // x=169, y=47
        pixel_data[47][170] = 4'b0111; // x=170, y=47
        pixel_data[47][171] = 4'b0111; // x=171, y=47
        pixel_data[47][172] = 4'b0111; // x=172, y=47
        pixel_data[47][173] = 4'b0111; // x=173, y=47
        pixel_data[47][174] = 4'b0111; // x=174, y=47
        pixel_data[47][175] = 4'b0111; // x=175, y=47
        pixel_data[47][176] = 4'b0111; // x=176, y=47
        pixel_data[47][177] = 4'b0111; // x=177, y=47
        pixel_data[47][178] = 4'b0111; // x=178, y=47
        pixel_data[47][179] = 4'b0111; // x=179, y=47
        pixel_data[48][0] = 4'b0111; // x=0, y=48
        pixel_data[48][1] = 4'b0111; // x=1, y=48
        pixel_data[48][2] = 4'b0111; // x=2, y=48
        pixel_data[48][3] = 4'b0111; // x=3, y=48
        pixel_data[48][4] = 4'b0111; // x=4, y=48
        pixel_data[48][5] = 4'b0111; // x=5, y=48
        pixel_data[48][6] = 4'b0111; // x=6, y=48
        pixel_data[48][7] = 4'b0111; // x=7, y=48
        pixel_data[48][8] = 4'b0111; // x=8, y=48
        pixel_data[48][9] = 4'b0111; // x=9, y=48
        pixel_data[48][10] = 4'b0111; // x=10, y=48
        pixel_data[48][11] = 4'b0111; // x=11, y=48
        pixel_data[48][12] = 4'b0111; // x=12, y=48
        pixel_data[48][13] = 4'b0111; // x=13, y=48
        pixel_data[48][14] = 4'b0111; // x=14, y=48
        pixel_data[48][15] = 4'b0111; // x=15, y=48
        pixel_data[48][16] = 4'b0111; // x=16, y=48
        pixel_data[48][17] = 4'b0111; // x=17, y=48
        pixel_data[48][18] = 4'b0111; // x=18, y=48
        pixel_data[48][19] = 4'b0111; // x=19, y=48
        pixel_data[48][20] = 4'b0111; // x=20, y=48
        pixel_data[48][21] = 4'b0111; // x=21, y=48
        pixel_data[48][22] = 4'b0111; // x=22, y=48
        pixel_data[48][23] = 4'b0111; // x=23, y=48
        pixel_data[48][24] = 4'b0111; // x=24, y=48
        pixel_data[48][25] = 4'b0111; // x=25, y=48
        pixel_data[48][26] = 4'b0111; // x=26, y=48
        pixel_data[48][27] = 4'b0111; // x=27, y=48
        pixel_data[48][28] = 4'b0111; // x=28, y=48
        pixel_data[48][29] = 4'b0111; // x=29, y=48
        pixel_data[48][30] = 4'b0111; // x=30, y=48
        pixel_data[48][31] = 4'b0111; // x=31, y=48
        pixel_data[48][32] = 4'b0111; // x=32, y=48
        pixel_data[48][33] = 4'b0111; // x=33, y=48
        pixel_data[48][34] = 4'b0111; // x=34, y=48
        pixel_data[48][35] = 4'b0111; // x=35, y=48
        pixel_data[48][36] = 4'b0111; // x=36, y=48
        pixel_data[48][37] = 4'b0111; // x=37, y=48
        pixel_data[48][38] = 4'b0111; // x=38, y=48
        pixel_data[48][39] = 4'b0111; // x=39, y=48
        pixel_data[48][40] = 4'b0111; // x=40, y=48
        pixel_data[48][41] = 4'b0111; // x=41, y=48
        pixel_data[48][42] = 4'b0111; // x=42, y=48
        pixel_data[48][43] = 4'b0111; // x=43, y=48
        pixel_data[48][44] = 4'b0111; // x=44, y=48
        pixel_data[48][45] = 4'b0111; // x=45, y=48
        pixel_data[48][46] = 4'b0111; // x=46, y=48
        pixel_data[48][47] = 4'b0111; // x=47, y=48
        pixel_data[48][48] = 4'b0111; // x=48, y=48
        pixel_data[48][49] = 4'b0111; // x=49, y=48
        pixel_data[48][50] = 4'b0111; // x=50, y=48
        pixel_data[48][51] = 4'b0111; // x=51, y=48
        pixel_data[48][52] = 4'b0111; // x=52, y=48
        pixel_data[48][53] = 4'b0111; // x=53, y=48
        pixel_data[48][54] = 4'b0111; // x=54, y=48
        pixel_data[48][55] = 4'b0111; // x=55, y=48
        pixel_data[48][56] = 4'b0111; // x=56, y=48
        pixel_data[48][57] = 4'b0111; // x=57, y=48
        pixel_data[48][58] = 4'b0111; // x=58, y=48
        pixel_data[48][59] = 4'b0111; // x=59, y=48
        pixel_data[48][60] = 4'b0111; // x=60, y=48
        pixel_data[48][61] = 4'b0111; // x=61, y=48
        pixel_data[48][62] = 4'b0111; // x=62, y=48
        pixel_data[48][63] = 4'b0111; // x=63, y=48
        pixel_data[48][64] = 4'b0111; // x=64, y=48
        pixel_data[48][65] = 4'b0111; // x=65, y=48
        pixel_data[48][66] = 4'b0111; // x=66, y=48
        pixel_data[48][67] = 4'b0111; // x=67, y=48
        pixel_data[48][68] = 4'b0111; // x=68, y=48
        pixel_data[48][69] = 4'b0111; // x=69, y=48
        pixel_data[48][70] = 4'b0111; // x=70, y=48
        pixel_data[48][71] = 4'b0111; // x=71, y=48
        pixel_data[48][72] = 4'b0111; // x=72, y=48
        pixel_data[48][73] = 4'b0111; // x=73, y=48
        pixel_data[48][74] = 4'b0111; // x=74, y=48
        pixel_data[48][75] = 4'b0111; // x=75, y=48
        pixel_data[48][76] = 4'b0111; // x=76, y=48
        pixel_data[48][77] = 4'b0111; // x=77, y=48
        pixel_data[48][78] = 4'b0111; // x=78, y=48
        pixel_data[48][79] = 4'b0111; // x=79, y=48
        pixel_data[48][80] = 4'b0111; // x=80, y=48
        pixel_data[48][81] = 4'b0111; // x=81, y=48
        pixel_data[48][82] = 4'b0111; // x=82, y=48
        pixel_data[48][83] = 4'b0111; // x=83, y=48
        pixel_data[48][84] = 4'b0111; // x=84, y=48
        pixel_data[48][85] = 4'b0111; // x=85, y=48
        pixel_data[48][86] = 4'b0111; // x=86, y=48
        pixel_data[48][87] = 4'b0111; // x=87, y=48
        pixel_data[48][88] = 4'b0111; // x=88, y=48
        pixel_data[48][89] = 4'b0111; // x=89, y=48
        pixel_data[48][90] = 4'b0111; // x=90, y=48
        pixel_data[48][91] = 4'b0111; // x=91, y=48
        pixel_data[48][92] = 4'b0111; // x=92, y=48
        pixel_data[48][93] = 4'b0111; // x=93, y=48
        pixel_data[48][94] = 4'b0111; // x=94, y=48
        pixel_data[48][95] = 4'b0111; // x=95, y=48
        pixel_data[48][96] = 4'b0111; // x=96, y=48
        pixel_data[48][97] = 4'b0111; // x=97, y=48
        pixel_data[48][98] = 4'b0111; // x=98, y=48
        pixel_data[48][99] = 4'b0111; // x=99, y=48
        pixel_data[48][100] = 4'b0111; // x=100, y=48
        pixel_data[48][101] = 4'b0111; // x=101, y=48
        pixel_data[48][102] = 4'b0111; // x=102, y=48
        pixel_data[48][103] = 4'b0111; // x=103, y=48
        pixel_data[48][104] = 4'b0111; // x=104, y=48
        pixel_data[48][105] = 4'b0111; // x=105, y=48
        pixel_data[48][106] = 4'b0111; // x=106, y=48
        pixel_data[48][107] = 4'b0111; // x=107, y=48
        pixel_data[48][108] = 4'b0111; // x=108, y=48
        pixel_data[48][109] = 4'b0111; // x=109, y=48
        pixel_data[48][110] = 4'b0111; // x=110, y=48
        pixel_data[48][111] = 4'b0111; // x=111, y=48
        pixel_data[48][112] = 4'b0111; // x=112, y=48
        pixel_data[48][113] = 4'b0111; // x=113, y=48
        pixel_data[48][114] = 4'b0111; // x=114, y=48
        pixel_data[48][115] = 4'b0111; // x=115, y=48
        pixel_data[48][116] = 4'b0111; // x=116, y=48
        pixel_data[48][117] = 4'b0111; // x=117, y=48
        pixel_data[48][118] = 4'b0111; // x=118, y=48
        pixel_data[48][119] = 4'b0111; // x=119, y=48
        pixel_data[48][120] = 4'b0111; // x=120, y=48
        pixel_data[48][121] = 4'b0111; // x=121, y=48
        pixel_data[48][122] = 4'b0111; // x=122, y=48
        pixel_data[48][123] = 4'b0111; // x=123, y=48
        pixel_data[48][124] = 4'b0111; // x=124, y=48
        pixel_data[48][125] = 4'b0111; // x=125, y=48
        pixel_data[48][126] = 4'b0111; // x=126, y=48
        pixel_data[48][127] = 4'b0111; // x=127, y=48
        pixel_data[48][128] = 4'b0111; // x=128, y=48
        pixel_data[48][129] = 4'b0111; // x=129, y=48
        pixel_data[48][130] = 4'b0111; // x=130, y=48
        pixel_data[48][131] = 4'b0111; // x=131, y=48
        pixel_data[48][132] = 4'b0111; // x=132, y=48
        pixel_data[48][133] = 4'b0111; // x=133, y=48
        pixel_data[48][134] = 4'b0111; // x=134, y=48
        pixel_data[48][135] = 4'b0111; // x=135, y=48
        pixel_data[48][136] = 4'b0111; // x=136, y=48
        pixel_data[48][137] = 4'b0111; // x=137, y=48
        pixel_data[48][138] = 4'b0111; // x=138, y=48
        pixel_data[48][139] = 4'b0111; // x=139, y=48
        pixel_data[48][140] = 4'b0111; // x=140, y=48
        pixel_data[48][141] = 4'b0111; // x=141, y=48
        pixel_data[48][142] = 4'b0111; // x=142, y=48
        pixel_data[48][143] = 4'b0111; // x=143, y=48
        pixel_data[48][144] = 4'b0111; // x=144, y=48
        pixel_data[48][145] = 4'b0111; // x=145, y=48
        pixel_data[48][146] = 4'b0111; // x=146, y=48
        pixel_data[48][147] = 4'b0111; // x=147, y=48
        pixel_data[48][148] = 4'b0111; // x=148, y=48
        pixel_data[48][149] = 4'b0111; // x=149, y=48
        pixel_data[48][150] = 4'b0111; // x=150, y=48
        pixel_data[48][151] = 4'b0111; // x=151, y=48
        pixel_data[48][152] = 4'b0111; // x=152, y=48
        pixel_data[48][153] = 4'b0111; // x=153, y=48
        pixel_data[48][154] = 4'b0111; // x=154, y=48
        pixel_data[48][155] = 4'b0111; // x=155, y=48
        pixel_data[48][156] = 4'b0111; // x=156, y=48
        pixel_data[48][157] = 4'b0111; // x=157, y=48
        pixel_data[48][158] = 4'b0111; // x=158, y=48
        pixel_data[48][159] = 4'b0111; // x=159, y=48
        pixel_data[48][160] = 4'b0111; // x=160, y=48
        pixel_data[48][161] = 4'b0111; // x=161, y=48
        pixel_data[48][162] = 4'b0111; // x=162, y=48
        pixel_data[48][163] = 4'b0111; // x=163, y=48
        pixel_data[48][164] = 4'b0111; // x=164, y=48
        pixel_data[48][165] = 4'b0111; // x=165, y=48
        pixel_data[48][166] = 4'b0111; // x=166, y=48
        pixel_data[48][167] = 4'b0111; // x=167, y=48
        pixel_data[48][168] = 4'b0111; // x=168, y=48
        pixel_data[48][169] = 4'b0111; // x=169, y=48
        pixel_data[48][170] = 4'b0111; // x=170, y=48
        pixel_data[48][171] = 4'b0111; // x=171, y=48
        pixel_data[48][172] = 4'b0111; // x=172, y=48
        pixel_data[48][173] = 4'b0111; // x=173, y=48
        pixel_data[48][174] = 4'b0111; // x=174, y=48
        pixel_data[48][175] = 4'b0111; // x=175, y=48
        pixel_data[48][176] = 4'b0111; // x=176, y=48
        pixel_data[48][177] = 4'b0111; // x=177, y=48
        pixel_data[48][178] = 4'b0111; // x=178, y=48
        pixel_data[48][179] = 4'b0111; // x=179, y=48
        pixel_data[49][0] = 4'b0111; // x=0, y=49
        pixel_data[49][1] = 4'b0111; // x=1, y=49
        pixel_data[49][2] = 4'b0111; // x=2, y=49
        pixel_data[49][3] = 4'b0111; // x=3, y=49
        pixel_data[49][4] = 4'b0111; // x=4, y=49
        pixel_data[49][5] = 4'b0111; // x=5, y=49
        pixel_data[49][6] = 4'b0111; // x=6, y=49
        pixel_data[49][7] = 4'b0111; // x=7, y=49
        pixel_data[49][8] = 4'b0111; // x=8, y=49
        pixel_data[49][9] = 4'b0111; // x=9, y=49
        pixel_data[49][10] = 4'b0111; // x=10, y=49
        pixel_data[49][11] = 4'b0111; // x=11, y=49
        pixel_data[49][12] = 4'b0111; // x=12, y=49
        pixel_data[49][13] = 4'b0111; // x=13, y=49
        pixel_data[49][14] = 4'b0111; // x=14, y=49
        pixel_data[49][15] = 4'b0111; // x=15, y=49
        pixel_data[49][16] = 4'b0111; // x=16, y=49
        pixel_data[49][17] = 4'b0111; // x=17, y=49
        pixel_data[49][18] = 4'b0111; // x=18, y=49
        pixel_data[49][19] = 4'b0111; // x=19, y=49
        pixel_data[49][20] = 4'b0111; // x=20, y=49
        pixel_data[49][21] = 4'b0111; // x=21, y=49
        pixel_data[49][22] = 4'b0111; // x=22, y=49
        pixel_data[49][23] = 4'b0111; // x=23, y=49
        pixel_data[49][24] = 4'b0111; // x=24, y=49
        pixel_data[49][25] = 4'b0111; // x=25, y=49
        pixel_data[49][26] = 4'b0111; // x=26, y=49
        pixel_data[49][27] = 4'b0111; // x=27, y=49
        pixel_data[49][28] = 4'b0111; // x=28, y=49
        pixel_data[49][29] = 4'b0111; // x=29, y=49
        pixel_data[49][30] = 4'b0111; // x=30, y=49
        pixel_data[49][31] = 4'b0111; // x=31, y=49
        pixel_data[49][32] = 4'b0111; // x=32, y=49
        pixel_data[49][33] = 4'b0111; // x=33, y=49
        pixel_data[49][34] = 4'b0111; // x=34, y=49
        pixel_data[49][35] = 4'b0111; // x=35, y=49
        pixel_data[49][36] = 4'b0111; // x=36, y=49
        pixel_data[49][37] = 4'b0111; // x=37, y=49
        pixel_data[49][38] = 4'b0111; // x=38, y=49
        pixel_data[49][39] = 4'b0111; // x=39, y=49
        pixel_data[49][40] = 4'b0111; // x=40, y=49
        pixel_data[49][41] = 4'b0111; // x=41, y=49
        pixel_data[49][42] = 4'b0111; // x=42, y=49
        pixel_data[49][43] = 4'b0111; // x=43, y=49
        pixel_data[49][44] = 4'b0111; // x=44, y=49
        pixel_data[49][45] = 4'b0111; // x=45, y=49
        pixel_data[49][46] = 4'b0111; // x=46, y=49
        pixel_data[49][47] = 4'b0111; // x=47, y=49
        pixel_data[49][48] = 4'b0111; // x=48, y=49
        pixel_data[49][49] = 4'b0111; // x=49, y=49
        pixel_data[49][50] = 4'b0111; // x=50, y=49
        pixel_data[49][51] = 4'b0111; // x=51, y=49
        pixel_data[49][52] = 4'b0111; // x=52, y=49
        pixel_data[49][53] = 4'b0111; // x=53, y=49
        pixel_data[49][54] = 4'b0111; // x=54, y=49
        pixel_data[49][55] = 4'b0111; // x=55, y=49
        pixel_data[49][56] = 4'b0111; // x=56, y=49
        pixel_data[49][57] = 4'b0111; // x=57, y=49
        pixel_data[49][58] = 4'b0111; // x=58, y=49
        pixel_data[49][59] = 4'b0111; // x=59, y=49
        pixel_data[49][60] = 4'b0111; // x=60, y=49
        pixel_data[49][61] = 4'b0111; // x=61, y=49
        pixel_data[49][62] = 4'b0111; // x=62, y=49
        pixel_data[49][63] = 4'b0111; // x=63, y=49
        pixel_data[49][64] = 4'b0111; // x=64, y=49
        pixel_data[49][65] = 4'b0111; // x=65, y=49
        pixel_data[49][66] = 4'b0111; // x=66, y=49
        pixel_data[49][67] = 4'b0111; // x=67, y=49
        pixel_data[49][68] = 4'b0111; // x=68, y=49
        pixel_data[49][69] = 4'b0111; // x=69, y=49
        pixel_data[49][70] = 4'b0111; // x=70, y=49
        pixel_data[49][71] = 4'b0111; // x=71, y=49
        pixel_data[49][72] = 4'b0111; // x=72, y=49
        pixel_data[49][73] = 4'b0111; // x=73, y=49
        pixel_data[49][74] = 4'b0111; // x=74, y=49
        pixel_data[49][75] = 4'b0111; // x=75, y=49
        pixel_data[49][76] = 4'b0111; // x=76, y=49
        pixel_data[49][77] = 4'b0111; // x=77, y=49
        pixel_data[49][78] = 4'b0111; // x=78, y=49
        pixel_data[49][79] = 4'b0111; // x=79, y=49
        pixel_data[49][80] = 4'b0111; // x=80, y=49
        pixel_data[49][81] = 4'b0111; // x=81, y=49
        pixel_data[49][82] = 4'b0111; // x=82, y=49
        pixel_data[49][83] = 4'b0111; // x=83, y=49
        pixel_data[49][84] = 4'b0111; // x=84, y=49
        pixel_data[49][85] = 4'b0111; // x=85, y=49
        pixel_data[49][86] = 4'b0111; // x=86, y=49
        pixel_data[49][87] = 4'b0111; // x=87, y=49
        pixel_data[49][88] = 4'b0111; // x=88, y=49
        pixel_data[49][89] = 4'b0111; // x=89, y=49
        pixel_data[49][90] = 4'b0111; // x=90, y=49
        pixel_data[49][91] = 4'b0111; // x=91, y=49
        pixel_data[49][92] = 4'b0111; // x=92, y=49
        pixel_data[49][93] = 4'b0111; // x=93, y=49
        pixel_data[49][94] = 4'b0111; // x=94, y=49
        pixel_data[49][95] = 4'b0111; // x=95, y=49
        pixel_data[49][96] = 4'b0111; // x=96, y=49
        pixel_data[49][97] = 4'b0111; // x=97, y=49
        pixel_data[49][98] = 4'b0111; // x=98, y=49
        pixel_data[49][99] = 4'b0111; // x=99, y=49
        pixel_data[49][100] = 4'b0111; // x=100, y=49
        pixel_data[49][101] = 4'b0111; // x=101, y=49
        pixel_data[49][102] = 4'b0111; // x=102, y=49
        pixel_data[49][103] = 4'b0111; // x=103, y=49
        pixel_data[49][104] = 4'b0111; // x=104, y=49
        pixel_data[49][105] = 4'b0111; // x=105, y=49
        pixel_data[49][106] = 4'b0111; // x=106, y=49
        pixel_data[49][107] = 4'b0111; // x=107, y=49
        pixel_data[49][108] = 4'b0111; // x=108, y=49
        pixel_data[49][109] = 4'b0111; // x=109, y=49
        pixel_data[49][110] = 4'b0111; // x=110, y=49
        pixel_data[49][111] = 4'b0111; // x=111, y=49
        pixel_data[49][112] = 4'b0111; // x=112, y=49
        pixel_data[49][113] = 4'b0111; // x=113, y=49
        pixel_data[49][114] = 4'b0111; // x=114, y=49
        pixel_data[49][115] = 4'b0111; // x=115, y=49
        pixel_data[49][116] = 4'b0111; // x=116, y=49
        pixel_data[49][117] = 4'b0111; // x=117, y=49
        pixel_data[49][118] = 4'b0111; // x=118, y=49
        pixel_data[49][119] = 4'b0111; // x=119, y=49
        pixel_data[49][120] = 4'b0111; // x=120, y=49
        pixel_data[49][121] = 4'b0111; // x=121, y=49
        pixel_data[49][122] = 4'b0111; // x=122, y=49
        pixel_data[49][123] = 4'b0111; // x=123, y=49
        pixel_data[49][124] = 4'b0111; // x=124, y=49
        pixel_data[49][125] = 4'b0111; // x=125, y=49
        pixel_data[49][126] = 4'b0111; // x=126, y=49
        pixel_data[49][127] = 4'b0111; // x=127, y=49
        pixel_data[49][128] = 4'b0111; // x=128, y=49
        pixel_data[49][129] = 4'b0111; // x=129, y=49
        pixel_data[49][130] = 4'b0111; // x=130, y=49
        pixel_data[49][131] = 4'b0111; // x=131, y=49
        pixel_data[49][132] = 4'b0111; // x=132, y=49
        pixel_data[49][133] = 4'b0111; // x=133, y=49
        pixel_data[49][134] = 4'b0111; // x=134, y=49
        pixel_data[49][135] = 4'b0111; // x=135, y=49
        pixel_data[49][136] = 4'b0111; // x=136, y=49
        pixel_data[49][137] = 4'b0111; // x=137, y=49
        pixel_data[49][138] = 4'b0111; // x=138, y=49
        pixel_data[49][139] = 4'b0111; // x=139, y=49
        pixel_data[49][140] = 4'b0111; // x=140, y=49
        pixel_data[49][141] = 4'b0111; // x=141, y=49
        pixel_data[49][142] = 4'b0111; // x=142, y=49
        pixel_data[49][143] = 4'b0111; // x=143, y=49
        pixel_data[49][144] = 4'b0111; // x=144, y=49
        pixel_data[49][145] = 4'b0111; // x=145, y=49
        pixel_data[49][146] = 4'b0111; // x=146, y=49
        pixel_data[49][147] = 4'b0111; // x=147, y=49
        pixel_data[49][148] = 4'b0111; // x=148, y=49
        pixel_data[49][149] = 4'b0111; // x=149, y=49
        pixel_data[49][150] = 4'b0111; // x=150, y=49
        pixel_data[49][151] = 4'b0111; // x=151, y=49
        pixel_data[49][152] = 4'b0111; // x=152, y=49
        pixel_data[49][153] = 4'b0111; // x=153, y=49
        pixel_data[49][154] = 4'b0111; // x=154, y=49
        pixel_data[49][155] = 4'b0111; // x=155, y=49
        pixel_data[49][156] = 4'b0111; // x=156, y=49
        pixel_data[49][157] = 4'b0111; // x=157, y=49
        pixel_data[49][158] = 4'b0111; // x=158, y=49
        pixel_data[49][159] = 4'b0111; // x=159, y=49
        pixel_data[49][160] = 4'b0111; // x=160, y=49
        pixel_data[49][161] = 4'b0111; // x=161, y=49
        pixel_data[49][162] = 4'b0111; // x=162, y=49
        pixel_data[49][163] = 4'b0111; // x=163, y=49
        pixel_data[49][164] = 4'b0111; // x=164, y=49
        pixel_data[49][165] = 4'b0111; // x=165, y=49
        pixel_data[49][166] = 4'b0111; // x=166, y=49
        pixel_data[49][167] = 4'b0111; // x=167, y=49
        pixel_data[49][168] = 4'b0111; // x=168, y=49
        pixel_data[49][169] = 4'b0111; // x=169, y=49
        pixel_data[49][170] = 4'b0111; // x=170, y=49
        pixel_data[49][171] = 4'b0111; // x=171, y=49
        pixel_data[49][172] = 4'b0111; // x=172, y=49
        pixel_data[49][173] = 4'b0111; // x=173, y=49
        pixel_data[49][174] = 4'b0111; // x=174, y=49
        pixel_data[49][175] = 4'b0111; // x=175, y=49
        pixel_data[49][176] = 4'b0111; // x=176, y=49
        pixel_data[49][177] = 4'b0111; // x=177, y=49
        pixel_data[49][178] = 4'b0111; // x=178, y=49
        pixel_data[49][179] = 4'b0111; // x=179, y=49
        pixel_data[50][0] = 4'b0111; // x=0, y=50
        pixel_data[50][1] = 4'b0111; // x=1, y=50
        pixel_data[50][2] = 4'b0111; // x=2, y=50
        pixel_data[50][3] = 4'b0111; // x=3, y=50
        pixel_data[50][4] = 4'b0111; // x=4, y=50
        pixel_data[50][5] = 4'b0111; // x=5, y=50
        pixel_data[50][6] = 4'b0111; // x=6, y=50
        pixel_data[50][7] = 4'b0111; // x=7, y=50
        pixel_data[50][8] = 4'b0111; // x=8, y=50
        pixel_data[50][9] = 4'b0111; // x=9, y=50
        pixel_data[50][10] = 4'b0111; // x=10, y=50
        pixel_data[50][11] = 4'b0111; // x=11, y=50
        pixel_data[50][12] = 4'b0111; // x=12, y=50
        pixel_data[50][13] = 4'b0111; // x=13, y=50
        pixel_data[50][14] = 4'b0111; // x=14, y=50
        pixel_data[50][15] = 4'b0111; // x=15, y=50
        pixel_data[50][16] = 4'b0111; // x=16, y=50
        pixel_data[50][17] = 4'b0111; // x=17, y=50
        pixel_data[50][18] = 4'b0111; // x=18, y=50
        pixel_data[50][19] = 4'b0111; // x=19, y=50
        pixel_data[50][20] = 4'b0111; // x=20, y=50
        pixel_data[50][21] = 4'b0111; // x=21, y=50
        pixel_data[50][22] = 4'b0111; // x=22, y=50
        pixel_data[50][23] = 4'b0111; // x=23, y=50
        pixel_data[50][24] = 4'b0111; // x=24, y=50
        pixel_data[50][25] = 4'b0111; // x=25, y=50
        pixel_data[50][26] = 4'b0111; // x=26, y=50
        pixel_data[50][27] = 4'b0111; // x=27, y=50
        pixel_data[50][28] = 4'b0111; // x=28, y=50
        pixel_data[50][29] = 4'b0111; // x=29, y=50
        pixel_data[50][30] = 4'b0111; // x=30, y=50
        pixel_data[50][31] = 4'b0111; // x=31, y=50
        pixel_data[50][32] = 4'b0111; // x=32, y=50
        pixel_data[50][33] = 4'b0111; // x=33, y=50
        pixel_data[50][34] = 4'b0111; // x=34, y=50
        pixel_data[50][35] = 4'b0111; // x=35, y=50
        pixel_data[50][36] = 4'b0111; // x=36, y=50
        pixel_data[50][37] = 4'b0111; // x=37, y=50
        pixel_data[50][38] = 4'b0111; // x=38, y=50
        pixel_data[50][39] = 4'b0111; // x=39, y=50
        pixel_data[50][40] = 4'b0111; // x=40, y=50
        pixel_data[50][41] = 4'b0111; // x=41, y=50
        pixel_data[50][42] = 4'b0111; // x=42, y=50
        pixel_data[50][43] = 4'b0111; // x=43, y=50
        pixel_data[50][44] = 4'b0111; // x=44, y=50
        pixel_data[50][45] = 4'b0111; // x=45, y=50
        pixel_data[50][46] = 4'b0111; // x=46, y=50
        pixel_data[50][47] = 4'b0111; // x=47, y=50
        pixel_data[50][48] = 4'b0111; // x=48, y=50
        pixel_data[50][49] = 4'b0111; // x=49, y=50
        pixel_data[50][50] = 4'b0111; // x=50, y=50
        pixel_data[50][51] = 4'b0111; // x=51, y=50
        pixel_data[50][52] = 4'b0111; // x=52, y=50
        pixel_data[50][53] = 4'b0111; // x=53, y=50
        pixel_data[50][54] = 4'b0111; // x=54, y=50
        pixel_data[50][55] = 4'b0111; // x=55, y=50
        pixel_data[50][56] = 4'b0111; // x=56, y=50
        pixel_data[50][57] = 4'b0111; // x=57, y=50
        pixel_data[50][58] = 4'b0111; // x=58, y=50
        pixel_data[50][59] = 4'b0111; // x=59, y=50
        pixel_data[50][60] = 4'b0111; // x=60, y=50
        pixel_data[50][61] = 4'b0111; // x=61, y=50
        pixel_data[50][62] = 4'b0111; // x=62, y=50
        pixel_data[50][63] = 4'b0111; // x=63, y=50
        pixel_data[50][64] = 4'b0111; // x=64, y=50
        pixel_data[50][65] = 4'b0111; // x=65, y=50
        pixel_data[50][66] = 4'b0111; // x=66, y=50
        pixel_data[50][67] = 4'b0111; // x=67, y=50
        pixel_data[50][68] = 4'b0111; // x=68, y=50
        pixel_data[50][69] = 4'b0111; // x=69, y=50
        pixel_data[50][70] = 4'b0111; // x=70, y=50
        pixel_data[50][71] = 4'b0111; // x=71, y=50
        pixel_data[50][72] = 4'b0111; // x=72, y=50
        pixel_data[50][73] = 4'b0111; // x=73, y=50
        pixel_data[50][74] = 4'b0111; // x=74, y=50
        pixel_data[50][75] = 4'b0111; // x=75, y=50
        pixel_data[50][76] = 4'b0111; // x=76, y=50
        pixel_data[50][77] = 4'b0111; // x=77, y=50
        pixel_data[50][78] = 4'b0111; // x=78, y=50
        pixel_data[50][79] = 4'b0111; // x=79, y=50
        pixel_data[50][80] = 4'b0111; // x=80, y=50
        pixel_data[50][81] = 4'b0111; // x=81, y=50
        pixel_data[50][82] = 4'b0111; // x=82, y=50
        pixel_data[50][83] = 4'b0111; // x=83, y=50
        pixel_data[50][84] = 4'b0111; // x=84, y=50
        pixel_data[50][85] = 4'b0111; // x=85, y=50
        pixel_data[50][86] = 4'b0111; // x=86, y=50
        pixel_data[50][87] = 4'b0111; // x=87, y=50
        pixel_data[50][88] = 4'b0111; // x=88, y=50
        pixel_data[50][89] = 4'b0111; // x=89, y=50
        pixel_data[50][90] = 4'b0111; // x=90, y=50
        pixel_data[50][91] = 4'b0111; // x=91, y=50
        pixel_data[50][92] = 4'b0111; // x=92, y=50
        pixel_data[50][93] = 4'b0111; // x=93, y=50
        pixel_data[50][94] = 4'b0111; // x=94, y=50
        pixel_data[50][95] = 4'b0111; // x=95, y=50
        pixel_data[50][96] = 4'b0111; // x=96, y=50
        pixel_data[50][97] = 4'b0111; // x=97, y=50
        pixel_data[50][98] = 4'b0111; // x=98, y=50
        pixel_data[50][99] = 4'b0111; // x=99, y=50
        pixel_data[50][100] = 4'b0111; // x=100, y=50
        pixel_data[50][101] = 4'b0111; // x=101, y=50
        pixel_data[50][102] = 4'b0111; // x=102, y=50
        pixel_data[50][103] = 4'b0111; // x=103, y=50
        pixel_data[50][104] = 4'b0111; // x=104, y=50
        pixel_data[50][105] = 4'b0111; // x=105, y=50
        pixel_data[50][106] = 4'b0111; // x=106, y=50
        pixel_data[50][107] = 4'b0111; // x=107, y=50
        pixel_data[50][108] = 4'b0111; // x=108, y=50
        pixel_data[50][109] = 4'b0111; // x=109, y=50
        pixel_data[50][110] = 4'b0111; // x=110, y=50
        pixel_data[50][111] = 4'b0111; // x=111, y=50
        pixel_data[50][112] = 4'b0111; // x=112, y=50
        pixel_data[50][113] = 4'b0111; // x=113, y=50
        pixel_data[50][114] = 4'b0111; // x=114, y=50
        pixel_data[50][115] = 4'b0111; // x=115, y=50
        pixel_data[50][116] = 4'b0111; // x=116, y=50
        pixel_data[50][117] = 4'b0111; // x=117, y=50
        pixel_data[50][118] = 4'b0111; // x=118, y=50
        pixel_data[50][119] = 4'b0111; // x=119, y=50
        pixel_data[50][120] = 4'b0111; // x=120, y=50
        pixel_data[50][121] = 4'b0111; // x=121, y=50
        pixel_data[50][122] = 4'b0111; // x=122, y=50
        pixel_data[50][123] = 4'b0111; // x=123, y=50
        pixel_data[50][124] = 4'b0111; // x=124, y=50
        pixel_data[50][125] = 4'b0111; // x=125, y=50
        pixel_data[50][126] = 4'b0111; // x=126, y=50
        pixel_data[50][127] = 4'b0111; // x=127, y=50
        pixel_data[50][128] = 4'b0111; // x=128, y=50
        pixel_data[50][129] = 4'b0111; // x=129, y=50
        pixel_data[50][130] = 4'b0111; // x=130, y=50
        pixel_data[50][131] = 4'b0111; // x=131, y=50
        pixel_data[50][132] = 4'b0111; // x=132, y=50
        pixel_data[50][133] = 4'b0111; // x=133, y=50
        pixel_data[50][134] = 4'b0111; // x=134, y=50
        pixel_data[50][135] = 4'b0111; // x=135, y=50
        pixel_data[50][136] = 4'b0111; // x=136, y=50
        pixel_data[50][137] = 4'b0111; // x=137, y=50
        pixel_data[50][138] = 4'b0111; // x=138, y=50
        pixel_data[50][139] = 4'b0111; // x=139, y=50
        pixel_data[50][140] = 4'b0111; // x=140, y=50
        pixel_data[50][141] = 4'b0111; // x=141, y=50
        pixel_data[50][142] = 4'b0111; // x=142, y=50
        pixel_data[50][143] = 4'b0111; // x=143, y=50
        pixel_data[50][144] = 4'b0111; // x=144, y=50
        pixel_data[50][145] = 4'b0111; // x=145, y=50
        pixel_data[50][146] = 4'b0111; // x=146, y=50
        pixel_data[50][147] = 4'b0111; // x=147, y=50
        pixel_data[50][148] = 4'b0111; // x=148, y=50
        pixel_data[50][149] = 4'b0111; // x=149, y=50
        pixel_data[50][150] = 4'b0111; // x=150, y=50
        pixel_data[50][151] = 4'b0111; // x=151, y=50
        pixel_data[50][152] = 4'b0111; // x=152, y=50
        pixel_data[50][153] = 4'b0111; // x=153, y=50
        pixel_data[50][154] = 4'b0111; // x=154, y=50
        pixel_data[50][155] = 4'b0111; // x=155, y=50
        pixel_data[50][156] = 4'b0111; // x=156, y=50
        pixel_data[50][157] = 4'b0111; // x=157, y=50
        pixel_data[50][158] = 4'b0111; // x=158, y=50
        pixel_data[50][159] = 4'b0111; // x=159, y=50
        pixel_data[50][160] = 4'b0111; // x=160, y=50
        pixel_data[50][161] = 4'b0111; // x=161, y=50
        pixel_data[50][162] = 4'b0111; // x=162, y=50
        pixel_data[50][163] = 4'b0111; // x=163, y=50
        pixel_data[50][164] = 4'b0111; // x=164, y=50
        pixel_data[50][165] = 4'b0111; // x=165, y=50
        pixel_data[50][166] = 4'b0111; // x=166, y=50
        pixel_data[50][167] = 4'b0111; // x=167, y=50
        pixel_data[50][168] = 4'b0111; // x=168, y=50
        pixel_data[50][169] = 4'b0111; // x=169, y=50
        pixel_data[50][170] = 4'b0111; // x=170, y=50
        pixel_data[50][171] = 4'b0111; // x=171, y=50
        pixel_data[50][172] = 4'b0111; // x=172, y=50
        pixel_data[50][173] = 4'b0111; // x=173, y=50
        pixel_data[50][174] = 4'b0111; // x=174, y=50
        pixel_data[50][175] = 4'b0111; // x=175, y=50
        pixel_data[50][176] = 4'b0111; // x=176, y=50
        pixel_data[50][177] = 4'b0111; // x=177, y=50
        pixel_data[50][178] = 4'b0111; // x=178, y=50
        pixel_data[50][179] = 4'b0111; // x=179, y=50
        pixel_data[51][0] = 4'b0111; // x=0, y=51
        pixel_data[51][1] = 4'b0111; // x=1, y=51
        pixel_data[51][2] = 4'b0111; // x=2, y=51
        pixel_data[51][3] = 4'b0111; // x=3, y=51
        pixel_data[51][4] = 4'b0111; // x=4, y=51
        pixel_data[51][5] = 4'b0111; // x=5, y=51
        pixel_data[51][6] = 4'b0111; // x=6, y=51
        pixel_data[51][7] = 4'b0111; // x=7, y=51
        pixel_data[51][8] = 4'b0111; // x=8, y=51
        pixel_data[51][9] = 4'b0111; // x=9, y=51
        pixel_data[51][10] = 4'b0111; // x=10, y=51
        pixel_data[51][11] = 4'b0111; // x=11, y=51
        pixel_data[51][12] = 4'b0111; // x=12, y=51
        pixel_data[51][13] = 4'b0111; // x=13, y=51
        pixel_data[51][14] = 4'b0111; // x=14, y=51
        pixel_data[51][15] = 4'b0111; // x=15, y=51
        pixel_data[51][16] = 4'b0111; // x=16, y=51
        pixel_data[51][17] = 4'b0111; // x=17, y=51
        pixel_data[51][18] = 4'b0111; // x=18, y=51
        pixel_data[51][19] = 4'b0111; // x=19, y=51
        pixel_data[51][20] = 4'b0111; // x=20, y=51
        pixel_data[51][21] = 4'b0111; // x=21, y=51
        pixel_data[51][22] = 4'b0111; // x=22, y=51
        pixel_data[51][23] = 4'b0111; // x=23, y=51
        pixel_data[51][24] = 4'b0111; // x=24, y=51
        pixel_data[51][25] = 4'b0111; // x=25, y=51
        pixel_data[51][26] = 4'b0111; // x=26, y=51
        pixel_data[51][27] = 4'b0111; // x=27, y=51
        pixel_data[51][28] = 4'b0111; // x=28, y=51
        pixel_data[51][29] = 4'b0111; // x=29, y=51
        pixel_data[51][30] = 4'b0111; // x=30, y=51
        pixel_data[51][31] = 4'b0111; // x=31, y=51
        pixel_data[51][32] = 4'b0111; // x=32, y=51
        pixel_data[51][33] = 4'b0111; // x=33, y=51
        pixel_data[51][34] = 4'b0111; // x=34, y=51
        pixel_data[51][35] = 4'b0111; // x=35, y=51
        pixel_data[51][36] = 4'b0111; // x=36, y=51
        pixel_data[51][37] = 4'b0111; // x=37, y=51
        pixel_data[51][38] = 4'b0111; // x=38, y=51
        pixel_data[51][39] = 4'b0111; // x=39, y=51
        pixel_data[51][40] = 4'b0111; // x=40, y=51
        pixel_data[51][41] = 4'b0111; // x=41, y=51
        pixel_data[51][42] = 4'b0111; // x=42, y=51
        pixel_data[51][43] = 4'b0111; // x=43, y=51
        pixel_data[51][44] = 4'b0111; // x=44, y=51
        pixel_data[51][45] = 4'b0111; // x=45, y=51
        pixel_data[51][46] = 4'b0111; // x=46, y=51
        pixel_data[51][47] = 4'b0111; // x=47, y=51
        pixel_data[51][48] = 4'b0111; // x=48, y=51
        pixel_data[51][49] = 4'b0111; // x=49, y=51
        pixel_data[51][50] = 4'b0111; // x=50, y=51
        pixel_data[51][51] = 4'b0111; // x=51, y=51
        pixel_data[51][52] = 4'b0111; // x=52, y=51
        pixel_data[51][53] = 4'b0111; // x=53, y=51
        pixel_data[51][54] = 4'b0111; // x=54, y=51
        pixel_data[51][55] = 4'b0111; // x=55, y=51
        pixel_data[51][56] = 4'b0111; // x=56, y=51
        pixel_data[51][57] = 4'b0111; // x=57, y=51
        pixel_data[51][58] = 4'b0111; // x=58, y=51
        pixel_data[51][59] = 4'b0111; // x=59, y=51
        pixel_data[51][60] = 4'b0111; // x=60, y=51
        pixel_data[51][61] = 4'b0111; // x=61, y=51
        pixel_data[51][62] = 4'b0111; // x=62, y=51
        pixel_data[51][63] = 4'b0111; // x=63, y=51
        pixel_data[51][64] = 4'b0111; // x=64, y=51
        pixel_data[51][65] = 4'b0111; // x=65, y=51
        pixel_data[51][66] = 4'b0111; // x=66, y=51
        pixel_data[51][67] = 4'b0111; // x=67, y=51
        pixel_data[51][68] = 4'b0111; // x=68, y=51
        pixel_data[51][69] = 4'b0111; // x=69, y=51
        pixel_data[51][70] = 4'b0111; // x=70, y=51
        pixel_data[51][71] = 4'b0111; // x=71, y=51
        pixel_data[51][72] = 4'b0111; // x=72, y=51
        pixel_data[51][73] = 4'b0111; // x=73, y=51
        pixel_data[51][74] = 4'b0111; // x=74, y=51
        pixel_data[51][75] = 4'b0111; // x=75, y=51
        pixel_data[51][76] = 4'b0111; // x=76, y=51
        pixel_data[51][77] = 4'b0111; // x=77, y=51
        pixel_data[51][78] = 4'b0111; // x=78, y=51
        pixel_data[51][79] = 4'b0111; // x=79, y=51
        pixel_data[51][80] = 4'b0111; // x=80, y=51
        pixel_data[51][81] = 4'b0111; // x=81, y=51
        pixel_data[51][82] = 4'b0111; // x=82, y=51
        pixel_data[51][83] = 4'b0111; // x=83, y=51
        pixel_data[51][84] = 4'b0111; // x=84, y=51
        pixel_data[51][85] = 4'b0111; // x=85, y=51
        pixel_data[51][86] = 4'b0111; // x=86, y=51
        pixel_data[51][87] = 4'b0111; // x=87, y=51
        pixel_data[51][88] = 4'b0111; // x=88, y=51
        pixel_data[51][89] = 4'b0111; // x=89, y=51
        pixel_data[51][90] = 4'b0111; // x=90, y=51
        pixel_data[51][91] = 4'b0111; // x=91, y=51
        pixel_data[51][92] = 4'b0111; // x=92, y=51
        pixel_data[51][93] = 4'b0111; // x=93, y=51
        pixel_data[51][94] = 4'b0111; // x=94, y=51
        pixel_data[51][95] = 4'b0111; // x=95, y=51
        pixel_data[51][96] = 4'b0111; // x=96, y=51
        pixel_data[51][97] = 4'b0111; // x=97, y=51
        pixel_data[51][98] = 4'b0111; // x=98, y=51
        pixel_data[51][99] = 4'b0111; // x=99, y=51
        pixel_data[51][100] = 4'b0111; // x=100, y=51
        pixel_data[51][101] = 4'b0111; // x=101, y=51
        pixel_data[51][102] = 4'b0111; // x=102, y=51
        pixel_data[51][103] = 4'b0111; // x=103, y=51
        pixel_data[51][104] = 4'b0111; // x=104, y=51
        pixel_data[51][105] = 4'b0111; // x=105, y=51
        pixel_data[51][106] = 4'b0111; // x=106, y=51
        pixel_data[51][107] = 4'b0111; // x=107, y=51
        pixel_data[51][108] = 4'b0111; // x=108, y=51
        pixel_data[51][109] = 4'b0111; // x=109, y=51
        pixel_data[51][110] = 4'b0111; // x=110, y=51
        pixel_data[51][111] = 4'b0111; // x=111, y=51
        pixel_data[51][112] = 4'b0111; // x=112, y=51
        pixel_data[51][113] = 4'b0111; // x=113, y=51
        pixel_data[51][114] = 4'b0111; // x=114, y=51
        pixel_data[51][115] = 4'b0111; // x=115, y=51
        pixel_data[51][116] = 4'b0111; // x=116, y=51
        pixel_data[51][117] = 4'b0111; // x=117, y=51
        pixel_data[51][118] = 4'b0111; // x=118, y=51
        pixel_data[51][119] = 4'b0111; // x=119, y=51
        pixel_data[51][120] = 4'b0111; // x=120, y=51
        pixel_data[51][121] = 4'b0111; // x=121, y=51
        pixel_data[51][122] = 4'b0111; // x=122, y=51
        pixel_data[51][123] = 4'b0111; // x=123, y=51
        pixel_data[51][124] = 4'b0111; // x=124, y=51
        pixel_data[51][125] = 4'b0111; // x=125, y=51
        pixel_data[51][126] = 4'b0111; // x=126, y=51
        pixel_data[51][127] = 4'b0111; // x=127, y=51
        pixel_data[51][128] = 4'b0111; // x=128, y=51
        pixel_data[51][129] = 4'b0111; // x=129, y=51
        pixel_data[51][130] = 4'b0111; // x=130, y=51
        pixel_data[51][131] = 4'b0111; // x=131, y=51
        pixel_data[51][132] = 4'b0111; // x=132, y=51
        pixel_data[51][133] = 4'b0111; // x=133, y=51
        pixel_data[51][134] = 4'b0111; // x=134, y=51
        pixel_data[51][135] = 4'b0111; // x=135, y=51
        pixel_data[51][136] = 4'b0111; // x=136, y=51
        pixel_data[51][137] = 4'b0111; // x=137, y=51
        pixel_data[51][138] = 4'b0111; // x=138, y=51
        pixel_data[51][139] = 4'b0111; // x=139, y=51
        pixel_data[51][140] = 4'b0111; // x=140, y=51
        pixel_data[51][141] = 4'b0111; // x=141, y=51
        pixel_data[51][142] = 4'b0111; // x=142, y=51
        pixel_data[51][143] = 4'b0111; // x=143, y=51
        pixel_data[51][144] = 4'b0111; // x=144, y=51
        pixel_data[51][145] = 4'b0111; // x=145, y=51
        pixel_data[51][146] = 4'b0111; // x=146, y=51
        pixel_data[51][147] = 4'b0111; // x=147, y=51
        pixel_data[51][148] = 4'b0111; // x=148, y=51
        pixel_data[51][149] = 4'b0111; // x=149, y=51
        pixel_data[51][150] = 4'b0111; // x=150, y=51
        pixel_data[51][151] = 4'b0111; // x=151, y=51
        pixel_data[51][152] = 4'b0111; // x=152, y=51
        pixel_data[51][153] = 4'b0111; // x=153, y=51
        pixel_data[51][154] = 4'b0111; // x=154, y=51
        pixel_data[51][155] = 4'b0111; // x=155, y=51
        pixel_data[51][156] = 4'b0111; // x=156, y=51
        pixel_data[51][157] = 4'b0111; // x=157, y=51
        pixel_data[51][158] = 4'b0111; // x=158, y=51
        pixel_data[51][159] = 4'b0111; // x=159, y=51
        pixel_data[51][160] = 4'b0111; // x=160, y=51
        pixel_data[51][161] = 4'b0111; // x=161, y=51
        pixel_data[51][162] = 4'b0111; // x=162, y=51
        pixel_data[51][163] = 4'b0111; // x=163, y=51
        pixel_data[51][164] = 4'b0111; // x=164, y=51
        pixel_data[51][165] = 4'b0111; // x=165, y=51
        pixel_data[51][166] = 4'b0111; // x=166, y=51
        pixel_data[51][167] = 4'b0111; // x=167, y=51
        pixel_data[51][168] = 4'b0111; // x=168, y=51
        pixel_data[51][169] = 4'b0111; // x=169, y=51
        pixel_data[51][170] = 4'b0111; // x=170, y=51
        pixel_data[51][171] = 4'b0111; // x=171, y=51
        pixel_data[51][172] = 4'b0111; // x=172, y=51
        pixel_data[51][173] = 4'b0111; // x=173, y=51
        pixel_data[51][174] = 4'b0111; // x=174, y=51
        pixel_data[51][175] = 4'b0111; // x=175, y=51
        pixel_data[51][176] = 4'b0111; // x=176, y=51
        pixel_data[51][177] = 4'b0111; // x=177, y=51
        pixel_data[51][178] = 4'b0111; // x=178, y=51
        pixel_data[51][179] = 4'b0111; // x=179, y=51
        pixel_data[52][0] = 4'b0111; // x=0, y=52
        pixel_data[52][1] = 4'b0111; // x=1, y=52
        pixel_data[52][2] = 4'b0111; // x=2, y=52
        pixel_data[52][3] = 4'b0111; // x=3, y=52
        pixel_data[52][4] = 4'b0111; // x=4, y=52
        pixel_data[52][5] = 4'b0111; // x=5, y=52
        pixel_data[52][6] = 4'b0111; // x=6, y=52
        pixel_data[52][7] = 4'b0111; // x=7, y=52
        pixel_data[52][8] = 4'b0111; // x=8, y=52
        pixel_data[52][9] = 4'b0111; // x=9, y=52
        pixel_data[52][10] = 4'b0111; // x=10, y=52
        pixel_data[52][11] = 4'b0111; // x=11, y=52
        pixel_data[52][12] = 4'b0111; // x=12, y=52
        pixel_data[52][13] = 4'b0111; // x=13, y=52
        pixel_data[52][14] = 4'b0111; // x=14, y=52
        pixel_data[52][15] = 4'b0111; // x=15, y=52
        pixel_data[52][16] = 4'b0111; // x=16, y=52
        pixel_data[52][17] = 4'b0111; // x=17, y=52
        pixel_data[52][18] = 4'b0111; // x=18, y=52
        pixel_data[52][19] = 4'b0111; // x=19, y=52
        pixel_data[52][20] = 4'b0111; // x=20, y=52
        pixel_data[52][21] = 4'b0111; // x=21, y=52
        pixel_data[52][22] = 4'b0111; // x=22, y=52
        pixel_data[52][23] = 4'b0111; // x=23, y=52
        pixel_data[52][24] = 4'b0111; // x=24, y=52
        pixel_data[52][25] = 4'b0111; // x=25, y=52
        pixel_data[52][26] = 4'b0111; // x=26, y=52
        pixel_data[52][27] = 4'b0111; // x=27, y=52
        pixel_data[52][28] = 4'b0111; // x=28, y=52
        pixel_data[52][29] = 4'b0111; // x=29, y=52
        pixel_data[52][30] = 4'b0111; // x=30, y=52
        pixel_data[52][31] = 4'b0111; // x=31, y=52
        pixel_data[52][32] = 4'b0111; // x=32, y=52
        pixel_data[52][33] = 4'b0111; // x=33, y=52
        pixel_data[52][34] = 4'b0111; // x=34, y=52
        pixel_data[52][35] = 4'b0111; // x=35, y=52
        pixel_data[52][36] = 4'b0111; // x=36, y=52
        pixel_data[52][37] = 4'b0111; // x=37, y=52
        pixel_data[52][38] = 4'b0111; // x=38, y=52
        pixel_data[52][39] = 4'b0111; // x=39, y=52
        pixel_data[52][40] = 4'b0111; // x=40, y=52
        pixel_data[52][41] = 4'b0111; // x=41, y=52
        pixel_data[52][42] = 4'b0111; // x=42, y=52
        pixel_data[52][43] = 4'b0111; // x=43, y=52
        pixel_data[52][44] = 4'b0111; // x=44, y=52
        pixel_data[52][45] = 4'b0111; // x=45, y=52
        pixel_data[52][46] = 4'b0111; // x=46, y=52
        pixel_data[52][47] = 4'b0111; // x=47, y=52
        pixel_data[52][48] = 4'b0111; // x=48, y=52
        pixel_data[52][49] = 4'b0111; // x=49, y=52
        pixel_data[52][50] = 4'b0111; // x=50, y=52
        pixel_data[52][51] = 4'b0111; // x=51, y=52
        pixel_data[52][52] = 4'b0111; // x=52, y=52
        pixel_data[52][53] = 4'b0111; // x=53, y=52
        pixel_data[52][54] = 4'b0111; // x=54, y=52
        pixel_data[52][55] = 4'b0111; // x=55, y=52
        pixel_data[52][56] = 4'b0111; // x=56, y=52
        pixel_data[52][57] = 4'b0111; // x=57, y=52
        pixel_data[52][58] = 4'b0111; // x=58, y=52
        pixel_data[52][59] = 4'b0111; // x=59, y=52
        pixel_data[52][60] = 4'b0111; // x=60, y=52
        pixel_data[52][61] = 4'b0111; // x=61, y=52
        pixel_data[52][62] = 4'b0111; // x=62, y=52
        pixel_data[52][63] = 4'b0111; // x=63, y=52
        pixel_data[52][64] = 4'b0111; // x=64, y=52
        pixel_data[52][65] = 4'b0111; // x=65, y=52
        pixel_data[52][66] = 4'b0111; // x=66, y=52
        pixel_data[52][67] = 4'b0111; // x=67, y=52
        pixel_data[52][68] = 4'b0111; // x=68, y=52
        pixel_data[52][69] = 4'b0111; // x=69, y=52
        pixel_data[52][70] = 4'b0111; // x=70, y=52
        pixel_data[52][71] = 4'b0111; // x=71, y=52
        pixel_data[52][72] = 4'b0111; // x=72, y=52
        pixel_data[52][73] = 4'b0111; // x=73, y=52
        pixel_data[52][74] = 4'b0111; // x=74, y=52
        pixel_data[52][75] = 4'b0111; // x=75, y=52
        pixel_data[52][76] = 4'b0111; // x=76, y=52
        pixel_data[52][77] = 4'b0111; // x=77, y=52
        pixel_data[52][78] = 4'b0111; // x=78, y=52
        pixel_data[52][79] = 4'b0111; // x=79, y=52
        pixel_data[52][80] = 4'b0111; // x=80, y=52
        pixel_data[52][81] = 4'b0111; // x=81, y=52
        pixel_data[52][82] = 4'b0111; // x=82, y=52
        pixel_data[52][83] = 4'b0111; // x=83, y=52
        pixel_data[52][84] = 4'b0111; // x=84, y=52
        pixel_data[52][85] = 4'b0111; // x=85, y=52
        pixel_data[52][86] = 4'b0111; // x=86, y=52
        pixel_data[52][87] = 4'b0111; // x=87, y=52
        pixel_data[52][88] = 4'b0111; // x=88, y=52
        pixel_data[52][89] = 4'b0111; // x=89, y=52
        pixel_data[52][90] = 4'b0111; // x=90, y=52
        pixel_data[52][91] = 4'b0111; // x=91, y=52
        pixel_data[52][92] = 4'b0111; // x=92, y=52
        pixel_data[52][93] = 4'b0111; // x=93, y=52
        pixel_data[52][94] = 4'b0111; // x=94, y=52
        pixel_data[52][95] = 4'b0111; // x=95, y=52
        pixel_data[52][96] = 4'b0111; // x=96, y=52
        pixel_data[52][97] = 4'b0111; // x=97, y=52
        pixel_data[52][98] = 4'b0111; // x=98, y=52
        pixel_data[52][99] = 4'b0111; // x=99, y=52
        pixel_data[52][100] = 4'b0111; // x=100, y=52
        pixel_data[52][101] = 4'b0111; // x=101, y=52
        pixel_data[52][102] = 4'b0111; // x=102, y=52
        pixel_data[52][103] = 4'b0111; // x=103, y=52
        pixel_data[52][104] = 4'b0111; // x=104, y=52
        pixel_data[52][105] = 4'b0111; // x=105, y=52
        pixel_data[52][106] = 4'b0111; // x=106, y=52
        pixel_data[52][107] = 4'b0111; // x=107, y=52
        pixel_data[52][108] = 4'b0111; // x=108, y=52
        pixel_data[52][109] = 4'b0111; // x=109, y=52
        pixel_data[52][110] = 4'b0111; // x=110, y=52
        pixel_data[52][111] = 4'b0111; // x=111, y=52
        pixel_data[52][112] = 4'b0111; // x=112, y=52
        pixel_data[52][113] = 4'b0111; // x=113, y=52
        pixel_data[52][114] = 4'b0111; // x=114, y=52
        pixel_data[52][115] = 4'b0111; // x=115, y=52
        pixel_data[52][116] = 4'b0111; // x=116, y=52
        pixel_data[52][117] = 4'b0111; // x=117, y=52
        pixel_data[52][118] = 4'b0111; // x=118, y=52
        pixel_data[52][119] = 4'b0111; // x=119, y=52
        pixel_data[52][120] = 4'b0111; // x=120, y=52
        pixel_data[52][121] = 4'b0111; // x=121, y=52
        pixel_data[52][122] = 4'b0111; // x=122, y=52
        pixel_data[52][123] = 4'b0111; // x=123, y=52
        pixel_data[52][124] = 4'b0111; // x=124, y=52
        pixel_data[52][125] = 4'b0111; // x=125, y=52
        pixel_data[52][126] = 4'b0111; // x=126, y=52
        pixel_data[52][127] = 4'b0111; // x=127, y=52
        pixel_data[52][128] = 4'b0111; // x=128, y=52
        pixel_data[52][129] = 4'b0111; // x=129, y=52
        pixel_data[52][130] = 4'b0111; // x=130, y=52
        pixel_data[52][131] = 4'b0111; // x=131, y=52
        pixel_data[52][132] = 4'b0111; // x=132, y=52
        pixel_data[52][133] = 4'b0111; // x=133, y=52
        pixel_data[52][134] = 4'b0111; // x=134, y=52
        pixel_data[52][135] = 4'b0111; // x=135, y=52
        pixel_data[52][136] = 4'b0111; // x=136, y=52
        pixel_data[52][137] = 4'b0111; // x=137, y=52
        pixel_data[52][138] = 4'b0111; // x=138, y=52
        pixel_data[52][139] = 4'b0111; // x=139, y=52
        pixel_data[52][140] = 4'b0111; // x=140, y=52
        pixel_data[52][141] = 4'b0111; // x=141, y=52
        pixel_data[52][142] = 4'b0111; // x=142, y=52
        pixel_data[52][143] = 4'b0111; // x=143, y=52
        pixel_data[52][144] = 4'b0111; // x=144, y=52
        pixel_data[52][145] = 4'b0111; // x=145, y=52
        pixel_data[52][146] = 4'b0111; // x=146, y=52
        pixel_data[52][147] = 4'b0111; // x=147, y=52
        pixel_data[52][148] = 4'b0111; // x=148, y=52
        pixel_data[52][149] = 4'b0111; // x=149, y=52
        pixel_data[52][150] = 4'b0111; // x=150, y=52
        pixel_data[52][151] = 4'b0111; // x=151, y=52
        pixel_data[52][152] = 4'b0111; // x=152, y=52
        pixel_data[52][153] = 4'b0111; // x=153, y=52
        pixel_data[52][154] = 4'b0111; // x=154, y=52
        pixel_data[52][155] = 4'b0111; // x=155, y=52
        pixel_data[52][156] = 4'b0111; // x=156, y=52
        pixel_data[52][157] = 4'b0111; // x=157, y=52
        pixel_data[52][158] = 4'b0111; // x=158, y=52
        pixel_data[52][159] = 4'b0111; // x=159, y=52
        pixel_data[52][160] = 4'b0111; // x=160, y=52
        pixel_data[52][161] = 4'b0111; // x=161, y=52
        pixel_data[52][162] = 4'b0111; // x=162, y=52
        pixel_data[52][163] = 4'b0111; // x=163, y=52
        pixel_data[52][164] = 4'b0111; // x=164, y=52
        pixel_data[52][165] = 4'b0111; // x=165, y=52
        pixel_data[52][166] = 4'b0111; // x=166, y=52
        pixel_data[52][167] = 4'b0111; // x=167, y=52
        pixel_data[52][168] = 4'b0111; // x=168, y=52
        pixel_data[52][169] = 4'b0111; // x=169, y=52
        pixel_data[52][170] = 4'b0111; // x=170, y=52
        pixel_data[52][171] = 4'b0111; // x=171, y=52
        pixel_data[52][172] = 4'b0111; // x=172, y=52
        pixel_data[52][173] = 4'b0111; // x=173, y=52
        pixel_data[52][174] = 4'b0111; // x=174, y=52
        pixel_data[52][175] = 4'b0111; // x=175, y=52
        pixel_data[52][176] = 4'b0111; // x=176, y=52
        pixel_data[52][177] = 4'b0111; // x=177, y=52
        pixel_data[52][178] = 4'b0111; // x=178, y=52
        pixel_data[52][179] = 4'b0111; // x=179, y=52
        pixel_data[53][0] = 4'b0111; // x=0, y=53
        pixel_data[53][1] = 4'b0111; // x=1, y=53
        pixel_data[53][2] = 4'b0111; // x=2, y=53
        pixel_data[53][3] = 4'b0111; // x=3, y=53
        pixel_data[53][4] = 4'b0111; // x=4, y=53
        pixel_data[53][5] = 4'b0111; // x=5, y=53
        pixel_data[53][6] = 4'b0111; // x=6, y=53
        pixel_data[53][7] = 4'b0111; // x=7, y=53
        pixel_data[53][8] = 4'b0111; // x=8, y=53
        pixel_data[53][9] = 4'b0111; // x=9, y=53
        pixel_data[53][10] = 4'b0111; // x=10, y=53
        pixel_data[53][11] = 4'b0111; // x=11, y=53
        pixel_data[53][12] = 4'b0111; // x=12, y=53
        pixel_data[53][13] = 4'b0111; // x=13, y=53
        pixel_data[53][14] = 4'b0111; // x=14, y=53
        pixel_data[53][15] = 4'b0111; // x=15, y=53
        pixel_data[53][16] = 4'b0111; // x=16, y=53
        pixel_data[53][17] = 4'b0111; // x=17, y=53
        pixel_data[53][18] = 4'b0111; // x=18, y=53
        pixel_data[53][19] = 4'b0111; // x=19, y=53
        pixel_data[53][20] = 4'b0111; // x=20, y=53
        pixel_data[53][21] = 4'b0111; // x=21, y=53
        pixel_data[53][22] = 4'b0111; // x=22, y=53
        pixel_data[53][23] = 4'b0111; // x=23, y=53
        pixel_data[53][24] = 4'b0111; // x=24, y=53
        pixel_data[53][25] = 4'b0111; // x=25, y=53
        pixel_data[53][26] = 4'b0111; // x=26, y=53
        pixel_data[53][27] = 4'b0111; // x=27, y=53
        pixel_data[53][28] = 4'b0111; // x=28, y=53
        pixel_data[53][29] = 4'b0111; // x=29, y=53
        pixel_data[53][30] = 4'b0111; // x=30, y=53
        pixel_data[53][31] = 4'b0111; // x=31, y=53
        pixel_data[53][32] = 4'b0111; // x=32, y=53
        pixel_data[53][33] = 4'b0111; // x=33, y=53
        pixel_data[53][34] = 4'b0111; // x=34, y=53
        pixel_data[53][35] = 4'b0111; // x=35, y=53
        pixel_data[53][36] = 4'b0111; // x=36, y=53
        pixel_data[53][37] = 4'b0111; // x=37, y=53
        pixel_data[53][38] = 4'b0111; // x=38, y=53
        pixel_data[53][39] = 4'b0111; // x=39, y=53
        pixel_data[53][40] = 4'b0111; // x=40, y=53
        pixel_data[53][41] = 4'b0111; // x=41, y=53
        pixel_data[53][42] = 4'b0111; // x=42, y=53
        pixel_data[53][43] = 4'b0111; // x=43, y=53
        pixel_data[53][44] = 4'b0111; // x=44, y=53
        pixel_data[53][45] = 4'b0111; // x=45, y=53
        pixel_data[53][46] = 4'b0111; // x=46, y=53
        pixel_data[53][47] = 4'b0111; // x=47, y=53
        pixel_data[53][48] = 4'b0111; // x=48, y=53
        pixel_data[53][49] = 4'b0111; // x=49, y=53
        pixel_data[53][50] = 4'b0111; // x=50, y=53
        pixel_data[53][51] = 4'b0111; // x=51, y=53
        pixel_data[53][52] = 4'b0111; // x=52, y=53
        pixel_data[53][53] = 4'b0111; // x=53, y=53
        pixel_data[53][54] = 4'b0111; // x=54, y=53
        pixel_data[53][55] = 4'b0111; // x=55, y=53
        pixel_data[53][56] = 4'b0111; // x=56, y=53
        pixel_data[53][57] = 4'b0111; // x=57, y=53
        pixel_data[53][58] = 4'b0111; // x=58, y=53
        pixel_data[53][59] = 4'b0111; // x=59, y=53
        pixel_data[53][60] = 4'b0111; // x=60, y=53
        pixel_data[53][61] = 4'b0111; // x=61, y=53
        pixel_data[53][62] = 4'b0111; // x=62, y=53
        pixel_data[53][63] = 4'b0111; // x=63, y=53
        pixel_data[53][64] = 4'b0111; // x=64, y=53
        pixel_data[53][65] = 4'b0111; // x=65, y=53
        pixel_data[53][66] = 4'b0111; // x=66, y=53
        pixel_data[53][67] = 4'b0111; // x=67, y=53
        pixel_data[53][68] = 4'b0111; // x=68, y=53
        pixel_data[53][69] = 4'b0111; // x=69, y=53
        pixel_data[53][70] = 4'b0111; // x=70, y=53
        pixel_data[53][71] = 4'b0111; // x=71, y=53
        pixel_data[53][72] = 4'b0111; // x=72, y=53
        pixel_data[53][73] = 4'b0111; // x=73, y=53
        pixel_data[53][74] = 4'b0111; // x=74, y=53
        pixel_data[53][75] = 4'b0111; // x=75, y=53
        pixel_data[53][76] = 4'b0111; // x=76, y=53
        pixel_data[53][77] = 4'b0111; // x=77, y=53
        pixel_data[53][78] = 4'b0111; // x=78, y=53
        pixel_data[53][79] = 4'b0111; // x=79, y=53
        pixel_data[53][80] = 4'b0111; // x=80, y=53
        pixel_data[53][81] = 4'b0111; // x=81, y=53
        pixel_data[53][82] = 4'b0111; // x=82, y=53
        pixel_data[53][83] = 4'b0111; // x=83, y=53
        pixel_data[53][84] = 4'b0111; // x=84, y=53
        pixel_data[53][85] = 4'b0111; // x=85, y=53
        pixel_data[53][86] = 4'b0111; // x=86, y=53
        pixel_data[53][87] = 4'b0111; // x=87, y=53
        pixel_data[53][88] = 4'b0111; // x=88, y=53
        pixel_data[53][89] = 4'b0111; // x=89, y=53
        pixel_data[53][90] = 4'b0111; // x=90, y=53
        pixel_data[53][91] = 4'b0111; // x=91, y=53
        pixel_data[53][92] = 4'b0111; // x=92, y=53
        pixel_data[53][93] = 4'b0111; // x=93, y=53
        pixel_data[53][94] = 4'b0111; // x=94, y=53
        pixel_data[53][95] = 4'b0111; // x=95, y=53
        pixel_data[53][96] = 4'b0111; // x=96, y=53
        pixel_data[53][97] = 4'b0111; // x=97, y=53
        pixel_data[53][98] = 4'b0111; // x=98, y=53
        pixel_data[53][99] = 4'b0111; // x=99, y=53
        pixel_data[53][100] = 4'b0111; // x=100, y=53
        pixel_data[53][101] = 4'b0111; // x=101, y=53
        pixel_data[53][102] = 4'b0111; // x=102, y=53
        pixel_data[53][103] = 4'b0111; // x=103, y=53
        pixel_data[53][104] = 4'b0111; // x=104, y=53
        pixel_data[53][105] = 4'b0111; // x=105, y=53
        pixel_data[53][106] = 4'b0111; // x=106, y=53
        pixel_data[53][107] = 4'b0111; // x=107, y=53
        pixel_data[53][108] = 4'b0111; // x=108, y=53
        pixel_data[53][109] = 4'b0111; // x=109, y=53
        pixel_data[53][110] = 4'b0111; // x=110, y=53
        pixel_data[53][111] = 4'b0111; // x=111, y=53
        pixel_data[53][112] = 4'b0111; // x=112, y=53
        pixel_data[53][113] = 4'b0111; // x=113, y=53
        pixel_data[53][114] = 4'b0111; // x=114, y=53
        pixel_data[53][115] = 4'b0111; // x=115, y=53
        pixel_data[53][116] = 4'b0111; // x=116, y=53
        pixel_data[53][117] = 4'b0111; // x=117, y=53
        pixel_data[53][118] = 4'b0111; // x=118, y=53
        pixel_data[53][119] = 4'b0111; // x=119, y=53
        pixel_data[53][120] = 4'b0111; // x=120, y=53
        pixel_data[53][121] = 4'b0111; // x=121, y=53
        pixel_data[53][122] = 4'b0111; // x=122, y=53
        pixel_data[53][123] = 4'b0111; // x=123, y=53
        pixel_data[53][124] = 4'b0111; // x=124, y=53
        pixel_data[53][125] = 4'b0111; // x=125, y=53
        pixel_data[53][126] = 4'b0111; // x=126, y=53
        pixel_data[53][127] = 4'b0111; // x=127, y=53
        pixel_data[53][128] = 4'b0111; // x=128, y=53
        pixel_data[53][129] = 4'b0111; // x=129, y=53
        pixel_data[53][130] = 4'b0111; // x=130, y=53
        pixel_data[53][131] = 4'b0111; // x=131, y=53
        pixel_data[53][132] = 4'b0111; // x=132, y=53
        pixel_data[53][133] = 4'b0111; // x=133, y=53
        pixel_data[53][134] = 4'b0111; // x=134, y=53
        pixel_data[53][135] = 4'b0111; // x=135, y=53
        pixel_data[53][136] = 4'b0111; // x=136, y=53
        pixel_data[53][137] = 4'b0111; // x=137, y=53
        pixel_data[53][138] = 4'b0111; // x=138, y=53
        pixel_data[53][139] = 4'b0111; // x=139, y=53
        pixel_data[53][140] = 4'b0111; // x=140, y=53
        pixel_data[53][141] = 4'b0111; // x=141, y=53
        pixel_data[53][142] = 4'b0111; // x=142, y=53
        pixel_data[53][143] = 4'b0111; // x=143, y=53
        pixel_data[53][144] = 4'b0111; // x=144, y=53
        pixel_data[53][145] = 4'b0111; // x=145, y=53
        pixel_data[53][146] = 4'b0111; // x=146, y=53
        pixel_data[53][147] = 4'b0111; // x=147, y=53
        pixel_data[53][148] = 4'b0111; // x=148, y=53
        pixel_data[53][149] = 4'b0111; // x=149, y=53
        pixel_data[53][150] = 4'b0111; // x=150, y=53
        pixel_data[53][151] = 4'b0111; // x=151, y=53
        pixel_data[53][152] = 4'b0111; // x=152, y=53
        pixel_data[53][153] = 4'b0111; // x=153, y=53
        pixel_data[53][154] = 4'b0111; // x=154, y=53
        pixel_data[53][155] = 4'b0111; // x=155, y=53
        pixel_data[53][156] = 4'b0111; // x=156, y=53
        pixel_data[53][157] = 4'b0111; // x=157, y=53
        pixel_data[53][158] = 4'b0111; // x=158, y=53
        pixel_data[53][159] = 4'b0111; // x=159, y=53
        pixel_data[53][160] = 4'b0111; // x=160, y=53
        pixel_data[53][161] = 4'b0111; // x=161, y=53
        pixel_data[53][162] = 4'b0111; // x=162, y=53
        pixel_data[53][163] = 4'b0111; // x=163, y=53
        pixel_data[53][164] = 4'b0111; // x=164, y=53
        pixel_data[53][165] = 4'b0111; // x=165, y=53
        pixel_data[53][166] = 4'b0111; // x=166, y=53
        pixel_data[53][167] = 4'b0111; // x=167, y=53
        pixel_data[53][168] = 4'b0111; // x=168, y=53
        pixel_data[53][169] = 4'b0111; // x=169, y=53
        pixel_data[53][170] = 4'b0111; // x=170, y=53
        pixel_data[53][171] = 4'b0111; // x=171, y=53
        pixel_data[53][172] = 4'b0111; // x=172, y=53
        pixel_data[53][173] = 4'b0111; // x=173, y=53
        pixel_data[53][174] = 4'b0111; // x=174, y=53
        pixel_data[53][175] = 4'b0111; // x=175, y=53
        pixel_data[53][176] = 4'b0111; // x=176, y=53
        pixel_data[53][177] = 4'b0111; // x=177, y=53
        pixel_data[53][178] = 4'b0111; // x=178, y=53
        pixel_data[53][179] = 4'b0111; // x=179, y=53
        pixel_data[54][0] = 4'b0111; // x=0, y=54
        pixel_data[54][1] = 4'b0111; // x=1, y=54
        pixel_data[54][2] = 4'b0111; // x=2, y=54
        pixel_data[54][3] = 4'b0111; // x=3, y=54
        pixel_data[54][4] = 4'b0111; // x=4, y=54
        pixel_data[54][5] = 4'b0111; // x=5, y=54
        pixel_data[54][6] = 4'b0111; // x=6, y=54
        pixel_data[54][7] = 4'b0111; // x=7, y=54
        pixel_data[54][8] = 4'b0111; // x=8, y=54
        pixel_data[54][9] = 4'b0111; // x=9, y=54
        pixel_data[54][10] = 4'b0111; // x=10, y=54
        pixel_data[54][11] = 4'b0111; // x=11, y=54
        pixel_data[54][12] = 4'b0111; // x=12, y=54
        pixel_data[54][13] = 4'b0111; // x=13, y=54
        pixel_data[54][14] = 4'b0111; // x=14, y=54
        pixel_data[54][15] = 4'b0111; // x=15, y=54
        pixel_data[54][16] = 4'b0111; // x=16, y=54
        pixel_data[54][17] = 4'b0111; // x=17, y=54
        pixel_data[54][18] = 4'b0111; // x=18, y=54
        pixel_data[54][19] = 4'b0111; // x=19, y=54
        pixel_data[54][20] = 4'b0111; // x=20, y=54
        pixel_data[54][21] = 4'b0111; // x=21, y=54
        pixel_data[54][22] = 4'b0111; // x=22, y=54
        pixel_data[54][23] = 4'b0111; // x=23, y=54
        pixel_data[54][24] = 4'b0111; // x=24, y=54
        pixel_data[54][25] = 4'b0111; // x=25, y=54
        pixel_data[54][26] = 4'b0111; // x=26, y=54
        pixel_data[54][27] = 4'b0111; // x=27, y=54
        pixel_data[54][28] = 4'b0111; // x=28, y=54
        pixel_data[54][29] = 4'b0111; // x=29, y=54
        pixel_data[54][30] = 4'b0111; // x=30, y=54
        pixel_data[54][31] = 4'b0111; // x=31, y=54
        pixel_data[54][32] = 4'b0111; // x=32, y=54
        pixel_data[54][33] = 4'b0111; // x=33, y=54
        pixel_data[54][34] = 4'b0111; // x=34, y=54
        pixel_data[54][35] = 4'b0111; // x=35, y=54
        pixel_data[54][36] = 4'b0111; // x=36, y=54
        pixel_data[54][37] = 4'b0111; // x=37, y=54
        pixel_data[54][38] = 4'b0111; // x=38, y=54
        pixel_data[54][39] = 4'b0111; // x=39, y=54
        pixel_data[54][40] = 4'b0111; // x=40, y=54
        pixel_data[54][41] = 4'b0111; // x=41, y=54
        pixel_data[54][42] = 4'b0111; // x=42, y=54
        pixel_data[54][43] = 4'b0111; // x=43, y=54
        pixel_data[54][44] = 4'b0111; // x=44, y=54
        pixel_data[54][45] = 4'b0111; // x=45, y=54
        pixel_data[54][46] = 4'b0111; // x=46, y=54
        pixel_data[54][47] = 4'b0111; // x=47, y=54
        pixel_data[54][48] = 4'b0111; // x=48, y=54
        pixel_data[54][49] = 4'b0111; // x=49, y=54
        pixel_data[54][50] = 4'b0111; // x=50, y=54
        pixel_data[54][51] = 4'b0111; // x=51, y=54
        pixel_data[54][52] = 4'b0111; // x=52, y=54
        pixel_data[54][53] = 4'b0111; // x=53, y=54
        pixel_data[54][54] = 4'b0111; // x=54, y=54
        pixel_data[54][55] = 4'b0111; // x=55, y=54
        pixel_data[54][56] = 4'b0111; // x=56, y=54
        pixel_data[54][57] = 4'b0111; // x=57, y=54
        pixel_data[54][58] = 4'b0111; // x=58, y=54
        pixel_data[54][59] = 4'b0111; // x=59, y=54
        pixel_data[54][60] = 4'b0111; // x=60, y=54
        pixel_data[54][61] = 4'b0111; // x=61, y=54
        pixel_data[54][62] = 4'b0111; // x=62, y=54
        pixel_data[54][63] = 4'b0111; // x=63, y=54
        pixel_data[54][64] = 4'b0111; // x=64, y=54
        pixel_data[54][65] = 4'b0111; // x=65, y=54
        pixel_data[54][66] = 4'b0111; // x=66, y=54
        pixel_data[54][67] = 4'b0111; // x=67, y=54
        pixel_data[54][68] = 4'b0111; // x=68, y=54
        pixel_data[54][69] = 4'b0111; // x=69, y=54
        pixel_data[54][70] = 4'b0111; // x=70, y=54
        pixel_data[54][71] = 4'b0111; // x=71, y=54
        pixel_data[54][72] = 4'b0111; // x=72, y=54
        pixel_data[54][73] = 4'b0111; // x=73, y=54
        pixel_data[54][74] = 4'b0111; // x=74, y=54
        pixel_data[54][75] = 4'b0111; // x=75, y=54
        pixel_data[54][76] = 4'b0111; // x=76, y=54
        pixel_data[54][77] = 4'b0111; // x=77, y=54
        pixel_data[54][78] = 4'b0111; // x=78, y=54
        pixel_data[54][79] = 4'b0111; // x=79, y=54
        pixel_data[54][80] = 4'b0111; // x=80, y=54
        pixel_data[54][81] = 4'b0111; // x=81, y=54
        pixel_data[54][82] = 4'b0111; // x=82, y=54
        pixel_data[54][83] = 4'b0111; // x=83, y=54
        pixel_data[54][84] = 4'b0111; // x=84, y=54
        pixel_data[54][85] = 4'b0111; // x=85, y=54
        pixel_data[54][86] = 4'b0111; // x=86, y=54
        pixel_data[54][87] = 4'b0111; // x=87, y=54
        pixel_data[54][88] = 4'b0111; // x=88, y=54
        pixel_data[54][89] = 4'b0111; // x=89, y=54
        pixel_data[54][90] = 4'b0111; // x=90, y=54
        pixel_data[54][91] = 4'b0111; // x=91, y=54
        pixel_data[54][92] = 4'b0111; // x=92, y=54
        pixel_data[54][93] = 4'b0111; // x=93, y=54
        pixel_data[54][94] = 4'b0111; // x=94, y=54
        pixel_data[54][95] = 4'b0111; // x=95, y=54
        pixel_data[54][96] = 4'b0111; // x=96, y=54
        pixel_data[54][97] = 4'b0111; // x=97, y=54
        pixel_data[54][98] = 4'b0111; // x=98, y=54
        pixel_data[54][99] = 4'b0111; // x=99, y=54
        pixel_data[54][100] = 4'b0111; // x=100, y=54
        pixel_data[54][101] = 4'b0111; // x=101, y=54
        pixel_data[54][102] = 4'b0111; // x=102, y=54
        pixel_data[54][103] = 4'b0111; // x=103, y=54
        pixel_data[54][104] = 4'b0111; // x=104, y=54
        pixel_data[54][105] = 4'b0111; // x=105, y=54
        pixel_data[54][106] = 4'b0111; // x=106, y=54
        pixel_data[54][107] = 4'b0111; // x=107, y=54
        pixel_data[54][108] = 4'b0111; // x=108, y=54
        pixel_data[54][109] = 4'b0111; // x=109, y=54
        pixel_data[54][110] = 4'b0111; // x=110, y=54
        pixel_data[54][111] = 4'b0111; // x=111, y=54
        pixel_data[54][112] = 4'b0111; // x=112, y=54
        pixel_data[54][113] = 4'b0111; // x=113, y=54
        pixel_data[54][114] = 4'b0111; // x=114, y=54
        pixel_data[54][115] = 4'b0111; // x=115, y=54
        pixel_data[54][116] = 4'b0111; // x=116, y=54
        pixel_data[54][117] = 4'b0111; // x=117, y=54
        pixel_data[54][118] = 4'b0111; // x=118, y=54
        pixel_data[54][119] = 4'b0111; // x=119, y=54
        pixel_data[54][120] = 4'b0111; // x=120, y=54
        pixel_data[54][121] = 4'b0111; // x=121, y=54
        pixel_data[54][122] = 4'b0111; // x=122, y=54
        pixel_data[54][123] = 4'b0111; // x=123, y=54
        pixel_data[54][124] = 4'b0111; // x=124, y=54
        pixel_data[54][125] = 4'b0111; // x=125, y=54
        pixel_data[54][126] = 4'b0111; // x=126, y=54
        pixel_data[54][127] = 4'b0111; // x=127, y=54
        pixel_data[54][128] = 4'b0111; // x=128, y=54
        pixel_data[54][129] = 4'b0111; // x=129, y=54
        pixel_data[54][130] = 4'b0111; // x=130, y=54
        pixel_data[54][131] = 4'b0111; // x=131, y=54
        pixel_data[54][132] = 4'b0111; // x=132, y=54
        pixel_data[54][133] = 4'b0111; // x=133, y=54
        pixel_data[54][134] = 4'b0111; // x=134, y=54
        pixel_data[54][135] = 4'b0111; // x=135, y=54
        pixel_data[54][136] = 4'b0111; // x=136, y=54
        pixel_data[54][137] = 4'b0111; // x=137, y=54
        pixel_data[54][138] = 4'b0111; // x=138, y=54
        pixel_data[54][139] = 4'b0111; // x=139, y=54
        pixel_data[54][140] = 4'b0111; // x=140, y=54
        pixel_data[54][141] = 4'b0111; // x=141, y=54
        pixel_data[54][142] = 4'b0111; // x=142, y=54
        pixel_data[54][143] = 4'b0111; // x=143, y=54
        pixel_data[54][144] = 4'b0111; // x=144, y=54
        pixel_data[54][145] = 4'b0111; // x=145, y=54
        pixel_data[54][146] = 4'b0111; // x=146, y=54
        pixel_data[54][147] = 4'b0111; // x=147, y=54
        pixel_data[54][148] = 4'b0111; // x=148, y=54
        pixel_data[54][149] = 4'b0111; // x=149, y=54
        pixel_data[54][150] = 4'b0111; // x=150, y=54
        pixel_data[54][151] = 4'b0111; // x=151, y=54
        pixel_data[54][152] = 4'b0111; // x=152, y=54
        pixel_data[54][153] = 4'b0111; // x=153, y=54
        pixel_data[54][154] = 4'b0111; // x=154, y=54
        pixel_data[54][155] = 4'b0111; // x=155, y=54
        pixel_data[54][156] = 4'b0111; // x=156, y=54
        pixel_data[54][157] = 4'b0111; // x=157, y=54
        pixel_data[54][158] = 4'b0111; // x=158, y=54
        pixel_data[54][159] = 4'b0111; // x=159, y=54
        pixel_data[54][160] = 4'b0111; // x=160, y=54
        pixel_data[54][161] = 4'b0111; // x=161, y=54
        pixel_data[54][162] = 4'b0111; // x=162, y=54
        pixel_data[54][163] = 4'b0111; // x=163, y=54
        pixel_data[54][164] = 4'b0111; // x=164, y=54
        pixel_data[54][165] = 4'b0111; // x=165, y=54
        pixel_data[54][166] = 4'b0111; // x=166, y=54
        pixel_data[54][167] = 4'b0111; // x=167, y=54
        pixel_data[54][168] = 4'b0111; // x=168, y=54
        pixel_data[54][169] = 4'b0111; // x=169, y=54
        pixel_data[54][170] = 4'b0111; // x=170, y=54
        pixel_data[54][171] = 4'b0111; // x=171, y=54
        pixel_data[54][172] = 4'b0111; // x=172, y=54
        pixel_data[54][173] = 4'b0111; // x=173, y=54
        pixel_data[54][174] = 4'b0111; // x=174, y=54
        pixel_data[54][175] = 4'b0111; // x=175, y=54
        pixel_data[54][176] = 4'b0111; // x=176, y=54
        pixel_data[54][177] = 4'b0111; // x=177, y=54
        pixel_data[54][178] = 4'b0111; // x=178, y=54
        pixel_data[54][179] = 4'b0111; // x=179, y=54
        pixel_data[55][0] = 4'b0111; // x=0, y=55
        pixel_data[55][1] = 4'b0111; // x=1, y=55
        pixel_data[55][2] = 4'b0111; // x=2, y=55
        pixel_data[55][3] = 4'b0111; // x=3, y=55
        pixel_data[55][4] = 4'b0111; // x=4, y=55
        pixel_data[55][5] = 4'b0111; // x=5, y=55
        pixel_data[55][6] = 4'b0111; // x=6, y=55
        pixel_data[55][7] = 4'b0111; // x=7, y=55
        pixel_data[55][8] = 4'b0111; // x=8, y=55
        pixel_data[55][9] = 4'b0111; // x=9, y=55
        pixel_data[55][10] = 4'b0111; // x=10, y=55
        pixel_data[55][11] = 4'b0111; // x=11, y=55
        pixel_data[55][12] = 4'b0111; // x=12, y=55
        pixel_data[55][13] = 4'b0111; // x=13, y=55
        pixel_data[55][14] = 4'b0111; // x=14, y=55
        pixel_data[55][15] = 4'b0111; // x=15, y=55
        pixel_data[55][16] = 4'b0111; // x=16, y=55
        pixel_data[55][17] = 4'b0111; // x=17, y=55
        pixel_data[55][18] = 4'b0111; // x=18, y=55
        pixel_data[55][19] = 4'b0111; // x=19, y=55
        pixel_data[55][20] = 4'b0111; // x=20, y=55
        pixel_data[55][21] = 4'b0111; // x=21, y=55
        pixel_data[55][22] = 4'b0111; // x=22, y=55
        pixel_data[55][23] = 4'b0111; // x=23, y=55
        pixel_data[55][24] = 4'b0111; // x=24, y=55
        pixel_data[55][25] = 4'b0111; // x=25, y=55
        pixel_data[55][26] = 4'b0111; // x=26, y=55
        pixel_data[55][27] = 4'b0111; // x=27, y=55
        pixel_data[55][28] = 4'b0111; // x=28, y=55
        pixel_data[55][29] = 4'b0111; // x=29, y=55
        pixel_data[55][30] = 4'b0111; // x=30, y=55
        pixel_data[55][31] = 4'b0111; // x=31, y=55
        pixel_data[55][32] = 4'b0111; // x=32, y=55
        pixel_data[55][33] = 4'b0111; // x=33, y=55
        pixel_data[55][34] = 4'b0111; // x=34, y=55
        pixel_data[55][35] = 4'b0111; // x=35, y=55
        pixel_data[55][36] = 4'b0111; // x=36, y=55
        pixel_data[55][37] = 4'b0111; // x=37, y=55
        pixel_data[55][38] = 4'b0111; // x=38, y=55
        pixel_data[55][39] = 4'b0111; // x=39, y=55
        pixel_data[55][40] = 4'b0111; // x=40, y=55
        pixel_data[55][41] = 4'b0111; // x=41, y=55
        pixel_data[55][42] = 4'b0111; // x=42, y=55
        pixel_data[55][43] = 4'b0111; // x=43, y=55
        pixel_data[55][44] = 4'b0111; // x=44, y=55
        pixel_data[55][45] = 4'b0111; // x=45, y=55
        pixel_data[55][46] = 4'b0111; // x=46, y=55
        pixel_data[55][47] = 4'b0111; // x=47, y=55
        pixel_data[55][48] = 4'b0111; // x=48, y=55
        pixel_data[55][49] = 4'b0111; // x=49, y=55
        pixel_data[55][50] = 4'b0111; // x=50, y=55
        pixel_data[55][51] = 4'b0111; // x=51, y=55
        pixel_data[55][52] = 4'b0111; // x=52, y=55
        pixel_data[55][53] = 4'b0111; // x=53, y=55
        pixel_data[55][54] = 4'b0111; // x=54, y=55
        pixel_data[55][55] = 4'b0111; // x=55, y=55
        pixel_data[55][56] = 4'b0111; // x=56, y=55
        pixel_data[55][57] = 4'b0111; // x=57, y=55
        pixel_data[55][58] = 4'b0111; // x=58, y=55
        pixel_data[55][59] = 4'b0111; // x=59, y=55
        pixel_data[55][60] = 4'b0111; // x=60, y=55
        pixel_data[55][61] = 4'b0111; // x=61, y=55
        pixel_data[55][62] = 4'b0111; // x=62, y=55
        pixel_data[55][63] = 4'b0111; // x=63, y=55
        pixel_data[55][64] = 4'b0111; // x=64, y=55
        pixel_data[55][65] = 4'b0111; // x=65, y=55
        pixel_data[55][66] = 4'b0111; // x=66, y=55
        pixel_data[55][67] = 4'b0111; // x=67, y=55
        pixel_data[55][68] = 4'b0111; // x=68, y=55
        pixel_data[55][69] = 4'b0111; // x=69, y=55
        pixel_data[55][70] = 4'b0111; // x=70, y=55
        pixel_data[55][71] = 4'b0111; // x=71, y=55
        pixel_data[55][72] = 4'b0111; // x=72, y=55
        pixel_data[55][73] = 4'b0111; // x=73, y=55
        pixel_data[55][74] = 4'b0111; // x=74, y=55
        pixel_data[55][75] = 4'b0111; // x=75, y=55
        pixel_data[55][76] = 4'b0111; // x=76, y=55
        pixel_data[55][77] = 4'b0111; // x=77, y=55
        pixel_data[55][78] = 4'b0111; // x=78, y=55
        pixel_data[55][79] = 4'b0111; // x=79, y=55
        pixel_data[55][80] = 4'b0111; // x=80, y=55
        pixel_data[55][81] = 4'b0111; // x=81, y=55
        pixel_data[55][82] = 4'b0111; // x=82, y=55
        pixel_data[55][83] = 4'b0111; // x=83, y=55
        pixel_data[55][84] = 4'b0111; // x=84, y=55
        pixel_data[55][85] = 4'b0111; // x=85, y=55
        pixel_data[55][86] = 4'b0111; // x=86, y=55
        pixel_data[55][87] = 4'b0111; // x=87, y=55
        pixel_data[55][88] = 4'b0111; // x=88, y=55
        pixel_data[55][89] = 4'b0111; // x=89, y=55
        pixel_data[55][90] = 4'b0111; // x=90, y=55
        pixel_data[55][91] = 4'b0111; // x=91, y=55
        pixel_data[55][92] = 4'b0111; // x=92, y=55
        pixel_data[55][93] = 4'b0111; // x=93, y=55
        pixel_data[55][94] = 4'b0111; // x=94, y=55
        pixel_data[55][95] = 4'b0111; // x=95, y=55
        pixel_data[55][96] = 4'b0111; // x=96, y=55
        pixel_data[55][97] = 4'b0111; // x=97, y=55
        pixel_data[55][98] = 4'b0111; // x=98, y=55
        pixel_data[55][99] = 4'b0111; // x=99, y=55
        pixel_data[55][100] = 4'b0111; // x=100, y=55
        pixel_data[55][101] = 4'b0111; // x=101, y=55
        pixel_data[55][102] = 4'b0111; // x=102, y=55
        pixel_data[55][103] = 4'b0111; // x=103, y=55
        pixel_data[55][104] = 4'b0111; // x=104, y=55
        pixel_data[55][105] = 4'b0111; // x=105, y=55
        pixel_data[55][106] = 4'b0111; // x=106, y=55
        pixel_data[55][107] = 4'b0111; // x=107, y=55
        pixel_data[55][108] = 4'b0111; // x=108, y=55
        pixel_data[55][109] = 4'b0111; // x=109, y=55
        pixel_data[55][110] = 4'b0111; // x=110, y=55
        pixel_data[55][111] = 4'b0111; // x=111, y=55
        pixel_data[55][112] = 4'b0111; // x=112, y=55
        pixel_data[55][113] = 4'b0111; // x=113, y=55
        pixel_data[55][114] = 4'b0111; // x=114, y=55
        pixel_data[55][115] = 4'b0111; // x=115, y=55
        pixel_data[55][116] = 4'b0111; // x=116, y=55
        pixel_data[55][117] = 4'b0111; // x=117, y=55
        pixel_data[55][118] = 4'b0111; // x=118, y=55
        pixel_data[55][119] = 4'b0111; // x=119, y=55
        pixel_data[55][120] = 4'b0111; // x=120, y=55
        pixel_data[55][121] = 4'b0111; // x=121, y=55
        pixel_data[55][122] = 4'b0111; // x=122, y=55
        pixel_data[55][123] = 4'b0111; // x=123, y=55
        pixel_data[55][124] = 4'b0111; // x=124, y=55
        pixel_data[55][125] = 4'b0111; // x=125, y=55
        pixel_data[55][126] = 4'b0111; // x=126, y=55
        pixel_data[55][127] = 4'b0111; // x=127, y=55
        pixel_data[55][128] = 4'b0111; // x=128, y=55
        pixel_data[55][129] = 4'b0111; // x=129, y=55
        pixel_data[55][130] = 4'b0111; // x=130, y=55
        pixel_data[55][131] = 4'b0111; // x=131, y=55
        pixel_data[55][132] = 4'b0111; // x=132, y=55
        pixel_data[55][133] = 4'b0111; // x=133, y=55
        pixel_data[55][134] = 4'b0111; // x=134, y=55
        pixel_data[55][135] = 4'b0111; // x=135, y=55
        pixel_data[55][136] = 4'b0111; // x=136, y=55
        pixel_data[55][137] = 4'b0111; // x=137, y=55
        pixel_data[55][138] = 4'b0111; // x=138, y=55
        pixel_data[55][139] = 4'b0111; // x=139, y=55
        pixel_data[55][140] = 4'b0111; // x=140, y=55
        pixel_data[55][141] = 4'b0111; // x=141, y=55
        pixel_data[55][142] = 4'b0111; // x=142, y=55
        pixel_data[55][143] = 4'b0111; // x=143, y=55
        pixel_data[55][144] = 4'b0111; // x=144, y=55
        pixel_data[55][145] = 4'b0111; // x=145, y=55
        pixel_data[55][146] = 4'b0111; // x=146, y=55
        pixel_data[55][147] = 4'b0111; // x=147, y=55
        pixel_data[55][148] = 4'b0111; // x=148, y=55
        pixel_data[55][149] = 4'b0111; // x=149, y=55
        pixel_data[55][150] = 4'b0111; // x=150, y=55
        pixel_data[55][151] = 4'b0111; // x=151, y=55
        pixel_data[55][152] = 4'b0111; // x=152, y=55
        pixel_data[55][153] = 4'b0111; // x=153, y=55
        pixel_data[55][154] = 4'b0111; // x=154, y=55
        pixel_data[55][155] = 4'b0111; // x=155, y=55
        pixel_data[55][156] = 4'b0111; // x=156, y=55
        pixel_data[55][157] = 4'b0111; // x=157, y=55
        pixel_data[55][158] = 4'b0111; // x=158, y=55
        pixel_data[55][159] = 4'b0111; // x=159, y=55
        pixel_data[55][160] = 4'b0111; // x=160, y=55
        pixel_data[55][161] = 4'b0111; // x=161, y=55
        pixel_data[55][162] = 4'b0111; // x=162, y=55
        pixel_data[55][163] = 4'b0111; // x=163, y=55
        pixel_data[55][164] = 4'b0111; // x=164, y=55
        pixel_data[55][165] = 4'b0111; // x=165, y=55
        pixel_data[55][166] = 4'b0111; // x=166, y=55
        pixel_data[55][167] = 4'b0111; // x=167, y=55
        pixel_data[55][168] = 4'b0111; // x=168, y=55
        pixel_data[55][169] = 4'b0111; // x=169, y=55
        pixel_data[55][170] = 4'b0111; // x=170, y=55
        pixel_data[55][171] = 4'b0111; // x=171, y=55
        pixel_data[55][172] = 4'b0111; // x=172, y=55
        pixel_data[55][173] = 4'b0111; // x=173, y=55
        pixel_data[55][174] = 4'b0111; // x=174, y=55
        pixel_data[55][175] = 4'b0111; // x=175, y=55
        pixel_data[55][176] = 4'b0111; // x=176, y=55
        pixel_data[55][177] = 4'b0111; // x=177, y=55
        pixel_data[55][178] = 4'b0111; // x=178, y=55
        pixel_data[55][179] = 4'b0111; // x=179, y=55
        pixel_data[56][0] = 4'b0111; // x=0, y=56
        pixel_data[56][1] = 4'b0111; // x=1, y=56
        pixel_data[56][2] = 4'b0111; // x=2, y=56
        pixel_data[56][3] = 4'b0111; // x=3, y=56
        pixel_data[56][4] = 4'b0111; // x=4, y=56
        pixel_data[56][5] = 4'b0111; // x=5, y=56
        pixel_data[56][6] = 4'b0111; // x=6, y=56
        pixel_data[56][7] = 4'b0111; // x=7, y=56
        pixel_data[56][8] = 4'b0111; // x=8, y=56
        pixel_data[56][9] = 4'b0111; // x=9, y=56
        pixel_data[56][10] = 4'b0111; // x=10, y=56
        pixel_data[56][11] = 4'b0111; // x=11, y=56
        pixel_data[56][12] = 4'b0111; // x=12, y=56
        pixel_data[56][13] = 4'b0111; // x=13, y=56
        pixel_data[56][14] = 4'b0111; // x=14, y=56
        pixel_data[56][15] = 4'b0111; // x=15, y=56
        pixel_data[56][16] = 4'b0111; // x=16, y=56
        pixel_data[56][17] = 4'b0111; // x=17, y=56
        pixel_data[56][18] = 4'b0111; // x=18, y=56
        pixel_data[56][19] = 4'b0111; // x=19, y=56
        pixel_data[56][20] = 4'b0111; // x=20, y=56
        pixel_data[56][21] = 4'b0111; // x=21, y=56
        pixel_data[56][22] = 4'b0111; // x=22, y=56
        pixel_data[56][23] = 4'b0111; // x=23, y=56
        pixel_data[56][24] = 4'b0111; // x=24, y=56
        pixel_data[56][25] = 4'b0111; // x=25, y=56
        pixel_data[56][26] = 4'b0111; // x=26, y=56
        pixel_data[56][27] = 4'b0111; // x=27, y=56
        pixel_data[56][28] = 4'b0111; // x=28, y=56
        pixel_data[56][29] = 4'b0111; // x=29, y=56
        pixel_data[56][30] = 4'b0111; // x=30, y=56
        pixel_data[56][31] = 4'b0111; // x=31, y=56
        pixel_data[56][32] = 4'b0111; // x=32, y=56
        pixel_data[56][33] = 4'b0111; // x=33, y=56
        pixel_data[56][34] = 4'b0111; // x=34, y=56
        pixel_data[56][35] = 4'b0111; // x=35, y=56
        pixel_data[56][36] = 4'b0111; // x=36, y=56
        pixel_data[56][37] = 4'b0111; // x=37, y=56
        pixel_data[56][38] = 4'b0111; // x=38, y=56
        pixel_data[56][39] = 4'b0111; // x=39, y=56
        pixel_data[56][40] = 4'b0111; // x=40, y=56
        pixel_data[56][41] = 4'b0111; // x=41, y=56
        pixel_data[56][42] = 4'b0111; // x=42, y=56
        pixel_data[56][43] = 4'b0111; // x=43, y=56
        pixel_data[56][44] = 4'b0111; // x=44, y=56
        pixel_data[56][45] = 4'b0111; // x=45, y=56
        pixel_data[56][46] = 4'b0111; // x=46, y=56
        pixel_data[56][47] = 4'b0111; // x=47, y=56
        pixel_data[56][48] = 4'b0111; // x=48, y=56
        pixel_data[56][49] = 4'b0111; // x=49, y=56
        pixel_data[56][50] = 4'b0111; // x=50, y=56
        pixel_data[56][51] = 4'b0111; // x=51, y=56
        pixel_data[56][52] = 4'b0111; // x=52, y=56
        pixel_data[56][53] = 4'b0111; // x=53, y=56
        pixel_data[56][54] = 4'b0111; // x=54, y=56
        pixel_data[56][55] = 4'b0111; // x=55, y=56
        pixel_data[56][56] = 4'b0111; // x=56, y=56
        pixel_data[56][57] = 4'b0111; // x=57, y=56
        pixel_data[56][58] = 4'b0111; // x=58, y=56
        pixel_data[56][59] = 4'b0111; // x=59, y=56
        pixel_data[56][60] = 4'b0111; // x=60, y=56
        pixel_data[56][61] = 4'b0111; // x=61, y=56
        pixel_data[56][62] = 4'b0111; // x=62, y=56
        pixel_data[56][63] = 4'b0111; // x=63, y=56
        pixel_data[56][64] = 4'b0111; // x=64, y=56
        pixel_data[56][65] = 4'b0111; // x=65, y=56
        pixel_data[56][66] = 4'b0111; // x=66, y=56
        pixel_data[56][67] = 4'b0111; // x=67, y=56
        pixel_data[56][68] = 4'b0111; // x=68, y=56
        pixel_data[56][69] = 4'b0111; // x=69, y=56
        pixel_data[56][70] = 4'b0111; // x=70, y=56
        pixel_data[56][71] = 4'b0111; // x=71, y=56
        pixel_data[56][72] = 4'b0111; // x=72, y=56
        pixel_data[56][73] = 4'b0111; // x=73, y=56
        pixel_data[56][74] = 4'b0111; // x=74, y=56
        pixel_data[56][75] = 4'b0111; // x=75, y=56
        pixel_data[56][76] = 4'b0111; // x=76, y=56
        pixel_data[56][77] = 4'b0111; // x=77, y=56
        pixel_data[56][78] = 4'b0111; // x=78, y=56
        pixel_data[56][79] = 4'b0111; // x=79, y=56
        pixel_data[56][80] = 4'b0111; // x=80, y=56
        pixel_data[56][81] = 4'b0111; // x=81, y=56
        pixel_data[56][82] = 4'b0111; // x=82, y=56
        pixel_data[56][83] = 4'b0111; // x=83, y=56
        pixel_data[56][84] = 4'b0111; // x=84, y=56
        pixel_data[56][85] = 4'b0111; // x=85, y=56
        pixel_data[56][86] = 4'b0111; // x=86, y=56
        pixel_data[56][87] = 4'b0111; // x=87, y=56
        pixel_data[56][88] = 4'b0111; // x=88, y=56
        pixel_data[56][89] = 4'b0111; // x=89, y=56
        pixel_data[56][90] = 4'b0111; // x=90, y=56
        pixel_data[56][91] = 4'b0111; // x=91, y=56
        pixel_data[56][92] = 4'b0111; // x=92, y=56
        pixel_data[56][93] = 4'b0111; // x=93, y=56
        pixel_data[56][94] = 4'b0111; // x=94, y=56
        pixel_data[56][95] = 4'b0111; // x=95, y=56
        pixel_data[56][96] = 4'b0111; // x=96, y=56
        pixel_data[56][97] = 4'b0111; // x=97, y=56
        pixel_data[56][98] = 4'b0111; // x=98, y=56
        pixel_data[56][99] = 4'b0111; // x=99, y=56
        pixel_data[56][100] = 4'b0111; // x=100, y=56
        pixel_data[56][101] = 4'b0111; // x=101, y=56
        pixel_data[56][102] = 4'b0111; // x=102, y=56
        pixel_data[56][103] = 4'b0111; // x=103, y=56
        pixel_data[56][104] = 4'b0111; // x=104, y=56
        pixel_data[56][105] = 4'b0111; // x=105, y=56
        pixel_data[56][106] = 4'b0111; // x=106, y=56
        pixel_data[56][107] = 4'b0111; // x=107, y=56
        pixel_data[56][108] = 4'b0111; // x=108, y=56
        pixel_data[56][109] = 4'b0111; // x=109, y=56
        pixel_data[56][110] = 4'b0111; // x=110, y=56
        pixel_data[56][111] = 4'b0111; // x=111, y=56
        pixel_data[56][112] = 4'b0111; // x=112, y=56
        pixel_data[56][113] = 4'b0111; // x=113, y=56
        pixel_data[56][114] = 4'b0111; // x=114, y=56
        pixel_data[56][115] = 4'b0111; // x=115, y=56
        pixel_data[56][116] = 4'b0111; // x=116, y=56
        pixel_data[56][117] = 4'b0111; // x=117, y=56
        pixel_data[56][118] = 4'b0111; // x=118, y=56
        pixel_data[56][119] = 4'b0111; // x=119, y=56
        pixel_data[56][120] = 4'b0111; // x=120, y=56
        pixel_data[56][121] = 4'b0111; // x=121, y=56
        pixel_data[56][122] = 4'b0111; // x=122, y=56
        pixel_data[56][123] = 4'b0111; // x=123, y=56
        pixel_data[56][124] = 4'b0111; // x=124, y=56
        pixel_data[56][125] = 4'b0111; // x=125, y=56
        pixel_data[56][126] = 4'b0111; // x=126, y=56
        pixel_data[56][127] = 4'b0111; // x=127, y=56
        pixel_data[56][128] = 4'b0111; // x=128, y=56
        pixel_data[56][129] = 4'b0111; // x=129, y=56
        pixel_data[56][130] = 4'b0111; // x=130, y=56
        pixel_data[56][131] = 4'b0111; // x=131, y=56
        pixel_data[56][132] = 4'b0111; // x=132, y=56
        pixel_data[56][133] = 4'b0111; // x=133, y=56
        pixel_data[56][134] = 4'b0111; // x=134, y=56
        pixel_data[56][135] = 4'b0111; // x=135, y=56
        pixel_data[56][136] = 4'b0111; // x=136, y=56
        pixel_data[56][137] = 4'b0111; // x=137, y=56
        pixel_data[56][138] = 4'b0111; // x=138, y=56
        pixel_data[56][139] = 4'b0111; // x=139, y=56
        pixel_data[56][140] = 4'b0111; // x=140, y=56
        pixel_data[56][141] = 4'b0111; // x=141, y=56
        pixel_data[56][142] = 4'b0111; // x=142, y=56
        pixel_data[56][143] = 4'b0111; // x=143, y=56
        pixel_data[56][144] = 4'b0111; // x=144, y=56
        pixel_data[56][145] = 4'b0111; // x=145, y=56
        pixel_data[56][146] = 4'b0111; // x=146, y=56
        pixel_data[56][147] = 4'b0111; // x=147, y=56
        pixel_data[56][148] = 4'b0111; // x=148, y=56
        pixel_data[56][149] = 4'b0111; // x=149, y=56
        pixel_data[56][150] = 4'b0111; // x=150, y=56
        pixel_data[56][151] = 4'b0111; // x=151, y=56
        pixel_data[56][152] = 4'b0111; // x=152, y=56
        pixel_data[56][153] = 4'b0111; // x=153, y=56
        pixel_data[56][154] = 4'b0111; // x=154, y=56
        pixel_data[56][155] = 4'b0111; // x=155, y=56
        pixel_data[56][156] = 4'b0111; // x=156, y=56
        pixel_data[56][157] = 4'b0111; // x=157, y=56
        pixel_data[56][158] = 4'b0111; // x=158, y=56
        pixel_data[56][159] = 4'b0111; // x=159, y=56
        pixel_data[56][160] = 4'b0111; // x=160, y=56
        pixel_data[56][161] = 4'b0111; // x=161, y=56
        pixel_data[56][162] = 4'b0111; // x=162, y=56
        pixel_data[56][163] = 4'b0111; // x=163, y=56
        pixel_data[56][164] = 4'b0111; // x=164, y=56
        pixel_data[56][165] = 4'b0111; // x=165, y=56
        pixel_data[56][166] = 4'b0111; // x=166, y=56
        pixel_data[56][167] = 4'b0111; // x=167, y=56
        pixel_data[56][168] = 4'b0111; // x=168, y=56
        pixel_data[56][169] = 4'b0111; // x=169, y=56
        pixel_data[56][170] = 4'b0111; // x=170, y=56
        pixel_data[56][171] = 4'b0111; // x=171, y=56
        pixel_data[56][172] = 4'b0111; // x=172, y=56
        pixel_data[56][173] = 4'b0111; // x=173, y=56
        pixel_data[56][174] = 4'b0111; // x=174, y=56
        pixel_data[56][175] = 4'b0111; // x=175, y=56
        pixel_data[56][176] = 4'b0111; // x=176, y=56
        pixel_data[56][177] = 4'b0111; // x=177, y=56
        pixel_data[56][178] = 4'b0111; // x=178, y=56
        pixel_data[56][179] = 4'b0111; // x=179, y=56
        pixel_data[57][0] = 4'b0111; // x=0, y=57
        pixel_data[57][1] = 4'b0111; // x=1, y=57
        pixel_data[57][2] = 4'b0111; // x=2, y=57
        pixel_data[57][3] = 4'b0111; // x=3, y=57
        pixel_data[57][4] = 4'b0111; // x=4, y=57
        pixel_data[57][5] = 4'b0111; // x=5, y=57
        pixel_data[57][6] = 4'b0111; // x=6, y=57
        pixel_data[57][7] = 4'b0111; // x=7, y=57
        pixel_data[57][8] = 4'b0111; // x=8, y=57
        pixel_data[57][9] = 4'b0111; // x=9, y=57
        pixel_data[57][10] = 4'b0111; // x=10, y=57
        pixel_data[57][11] = 4'b0111; // x=11, y=57
        pixel_data[57][12] = 4'b0111; // x=12, y=57
        pixel_data[57][13] = 4'b0111; // x=13, y=57
        pixel_data[57][14] = 4'b0111; // x=14, y=57
        pixel_data[57][15] = 4'b0111; // x=15, y=57
        pixel_data[57][16] = 4'b0111; // x=16, y=57
        pixel_data[57][17] = 4'b0111; // x=17, y=57
        pixel_data[57][18] = 4'b0111; // x=18, y=57
        pixel_data[57][19] = 4'b0111; // x=19, y=57
        pixel_data[57][20] = 4'b0111; // x=20, y=57
        pixel_data[57][21] = 4'b0111; // x=21, y=57
        pixel_data[57][22] = 4'b0111; // x=22, y=57
        pixel_data[57][23] = 4'b0111; // x=23, y=57
        pixel_data[57][24] = 4'b0111; // x=24, y=57
        pixel_data[57][25] = 4'b0111; // x=25, y=57
        pixel_data[57][26] = 4'b0111; // x=26, y=57
        pixel_data[57][27] = 4'b0111; // x=27, y=57
        pixel_data[57][28] = 4'b0111; // x=28, y=57
        pixel_data[57][29] = 4'b0111; // x=29, y=57
        pixel_data[57][30] = 4'b0111; // x=30, y=57
        pixel_data[57][31] = 4'b0111; // x=31, y=57
        pixel_data[57][32] = 4'b0111; // x=32, y=57
        pixel_data[57][33] = 4'b0111; // x=33, y=57
        pixel_data[57][34] = 4'b0111; // x=34, y=57
        pixel_data[57][35] = 4'b0111; // x=35, y=57
        pixel_data[57][36] = 4'b0111; // x=36, y=57
        pixel_data[57][37] = 4'b0111; // x=37, y=57
        pixel_data[57][38] = 4'b0111; // x=38, y=57
        pixel_data[57][39] = 4'b0111; // x=39, y=57
        pixel_data[57][40] = 4'b0111; // x=40, y=57
        pixel_data[57][41] = 4'b0111; // x=41, y=57
        pixel_data[57][42] = 4'b0111; // x=42, y=57
        pixel_data[57][43] = 4'b0111; // x=43, y=57
        pixel_data[57][44] = 4'b0111; // x=44, y=57
        pixel_data[57][45] = 4'b0111; // x=45, y=57
        pixel_data[57][46] = 4'b0111; // x=46, y=57
        pixel_data[57][47] = 4'b0111; // x=47, y=57
        pixel_data[57][48] = 4'b0111; // x=48, y=57
        pixel_data[57][49] = 4'b0111; // x=49, y=57
        pixel_data[57][50] = 4'b0111; // x=50, y=57
        pixel_data[57][51] = 4'b0111; // x=51, y=57
        pixel_data[57][52] = 4'b0111; // x=52, y=57
        pixel_data[57][53] = 4'b0111; // x=53, y=57
        pixel_data[57][54] = 4'b0111; // x=54, y=57
        pixel_data[57][55] = 4'b0111; // x=55, y=57
        pixel_data[57][56] = 4'b0111; // x=56, y=57
        pixel_data[57][57] = 4'b0111; // x=57, y=57
        pixel_data[57][58] = 4'b0111; // x=58, y=57
        pixel_data[57][59] = 4'b0111; // x=59, y=57
        pixel_data[57][60] = 4'b0111; // x=60, y=57
        pixel_data[57][61] = 4'b0111; // x=61, y=57
        pixel_data[57][62] = 4'b0111; // x=62, y=57
        pixel_data[57][63] = 4'b0111; // x=63, y=57
        pixel_data[57][64] = 4'b0111; // x=64, y=57
        pixel_data[57][65] = 4'b0111; // x=65, y=57
        pixel_data[57][66] = 4'b0111; // x=66, y=57
        pixel_data[57][67] = 4'b0111; // x=67, y=57
        pixel_data[57][68] = 4'b0111; // x=68, y=57
        pixel_data[57][69] = 4'b0111; // x=69, y=57
        pixel_data[57][70] = 4'b0111; // x=70, y=57
        pixel_data[57][71] = 4'b0111; // x=71, y=57
        pixel_data[57][72] = 4'b0111; // x=72, y=57
        pixel_data[57][73] = 4'b0111; // x=73, y=57
        pixel_data[57][74] = 4'b0111; // x=74, y=57
        pixel_data[57][75] = 4'b0111; // x=75, y=57
        pixel_data[57][76] = 4'b0111; // x=76, y=57
        pixel_data[57][77] = 4'b0111; // x=77, y=57
        pixel_data[57][78] = 4'b0111; // x=78, y=57
        pixel_data[57][79] = 4'b0111; // x=79, y=57
        pixel_data[57][80] = 4'b0111; // x=80, y=57
        pixel_data[57][81] = 4'b0111; // x=81, y=57
        pixel_data[57][82] = 4'b0111; // x=82, y=57
        pixel_data[57][83] = 4'b0111; // x=83, y=57
        pixel_data[57][84] = 4'b0111; // x=84, y=57
        pixel_data[57][85] = 4'b0111; // x=85, y=57
        pixel_data[57][86] = 4'b0111; // x=86, y=57
        pixel_data[57][87] = 4'b0111; // x=87, y=57
        pixel_data[57][88] = 4'b0111; // x=88, y=57
        pixel_data[57][89] = 4'b0111; // x=89, y=57
        pixel_data[57][90] = 4'b0111; // x=90, y=57
        pixel_data[57][91] = 4'b0111; // x=91, y=57
        pixel_data[57][92] = 4'b0111; // x=92, y=57
        pixel_data[57][93] = 4'b0111; // x=93, y=57
        pixel_data[57][94] = 4'b0111; // x=94, y=57
        pixel_data[57][95] = 4'b0111; // x=95, y=57
        pixel_data[57][96] = 4'b0111; // x=96, y=57
        pixel_data[57][97] = 4'b0111; // x=97, y=57
        pixel_data[57][98] = 4'b0111; // x=98, y=57
        pixel_data[57][99] = 4'b0111; // x=99, y=57
        pixel_data[57][100] = 4'b0111; // x=100, y=57
        pixel_data[57][101] = 4'b0111; // x=101, y=57
        pixel_data[57][102] = 4'b0111; // x=102, y=57
        pixel_data[57][103] = 4'b0111; // x=103, y=57
        pixel_data[57][104] = 4'b0111; // x=104, y=57
        pixel_data[57][105] = 4'b0111; // x=105, y=57
        pixel_data[57][106] = 4'b0111; // x=106, y=57
        pixel_data[57][107] = 4'b0111; // x=107, y=57
        pixel_data[57][108] = 4'b0111; // x=108, y=57
        pixel_data[57][109] = 4'b0111; // x=109, y=57
        pixel_data[57][110] = 4'b0111; // x=110, y=57
        pixel_data[57][111] = 4'b0111; // x=111, y=57
        pixel_data[57][112] = 4'b0111; // x=112, y=57
        pixel_data[57][113] = 4'b0111; // x=113, y=57
        pixel_data[57][114] = 4'b0111; // x=114, y=57
        pixel_data[57][115] = 4'b0111; // x=115, y=57
        pixel_data[57][116] = 4'b0111; // x=116, y=57
        pixel_data[57][117] = 4'b0111; // x=117, y=57
        pixel_data[57][118] = 4'b0111; // x=118, y=57
        pixel_data[57][119] = 4'b0111; // x=119, y=57
        pixel_data[57][120] = 4'b0111; // x=120, y=57
        pixel_data[57][121] = 4'b0111; // x=121, y=57
        pixel_data[57][122] = 4'b0111; // x=122, y=57
        pixel_data[57][123] = 4'b0111; // x=123, y=57
        pixel_data[57][124] = 4'b0111; // x=124, y=57
        pixel_data[57][125] = 4'b0111; // x=125, y=57
        pixel_data[57][126] = 4'b0111; // x=126, y=57
        pixel_data[57][127] = 4'b0111; // x=127, y=57
        pixel_data[57][128] = 4'b0111; // x=128, y=57
        pixel_data[57][129] = 4'b0111; // x=129, y=57
        pixel_data[57][130] = 4'b0111; // x=130, y=57
        pixel_data[57][131] = 4'b0111; // x=131, y=57
        pixel_data[57][132] = 4'b0111; // x=132, y=57
        pixel_data[57][133] = 4'b0111; // x=133, y=57
        pixel_data[57][134] = 4'b0111; // x=134, y=57
        pixel_data[57][135] = 4'b0111; // x=135, y=57
        pixel_data[57][136] = 4'b0111; // x=136, y=57
        pixel_data[57][137] = 4'b0111; // x=137, y=57
        pixel_data[57][138] = 4'b0111; // x=138, y=57
        pixel_data[57][139] = 4'b0111; // x=139, y=57
        pixel_data[57][140] = 4'b0111; // x=140, y=57
        pixel_data[57][141] = 4'b0111; // x=141, y=57
        pixel_data[57][142] = 4'b0111; // x=142, y=57
        pixel_data[57][143] = 4'b0111; // x=143, y=57
        pixel_data[57][144] = 4'b0111; // x=144, y=57
        pixel_data[57][145] = 4'b0111; // x=145, y=57
        pixel_data[57][146] = 4'b0111; // x=146, y=57
        pixel_data[57][147] = 4'b0111; // x=147, y=57
        pixel_data[57][148] = 4'b0111; // x=148, y=57
        pixel_data[57][149] = 4'b0111; // x=149, y=57
        pixel_data[57][150] = 4'b0111; // x=150, y=57
        pixel_data[57][151] = 4'b0111; // x=151, y=57
        pixel_data[57][152] = 4'b0111; // x=152, y=57
        pixel_data[57][153] = 4'b0111; // x=153, y=57
        pixel_data[57][154] = 4'b0111; // x=154, y=57
        pixel_data[57][155] = 4'b0111; // x=155, y=57
        pixel_data[57][156] = 4'b0111; // x=156, y=57
        pixel_data[57][157] = 4'b0111; // x=157, y=57
        pixel_data[57][158] = 4'b0111; // x=158, y=57
        pixel_data[57][159] = 4'b0111; // x=159, y=57
        pixel_data[57][160] = 4'b0111; // x=160, y=57
        pixel_data[57][161] = 4'b0111; // x=161, y=57
        pixel_data[57][162] = 4'b0111; // x=162, y=57
        pixel_data[57][163] = 4'b0111; // x=163, y=57
        pixel_data[57][164] = 4'b0111; // x=164, y=57
        pixel_data[57][165] = 4'b0111; // x=165, y=57
        pixel_data[57][166] = 4'b0111; // x=166, y=57
        pixel_data[57][167] = 4'b0111; // x=167, y=57
        pixel_data[57][168] = 4'b0111; // x=168, y=57
        pixel_data[57][169] = 4'b0111; // x=169, y=57
        pixel_data[57][170] = 4'b0111; // x=170, y=57
        pixel_data[57][171] = 4'b0111; // x=171, y=57
        pixel_data[57][172] = 4'b0111; // x=172, y=57
        pixel_data[57][173] = 4'b0111; // x=173, y=57
        pixel_data[57][174] = 4'b0111; // x=174, y=57
        pixel_data[57][175] = 4'b0111; // x=175, y=57
        pixel_data[57][176] = 4'b0111; // x=176, y=57
        pixel_data[57][177] = 4'b0111; // x=177, y=57
        pixel_data[57][178] = 4'b0111; // x=178, y=57
        pixel_data[57][179] = 4'b0111; // x=179, y=57
        pixel_data[58][0] = 4'b0111; // x=0, y=58
        pixel_data[58][1] = 4'b0111; // x=1, y=58
        pixel_data[58][2] = 4'b0111; // x=2, y=58
        pixel_data[58][3] = 4'b0111; // x=3, y=58
        pixel_data[58][4] = 4'b0111; // x=4, y=58
        pixel_data[58][5] = 4'b0111; // x=5, y=58
        pixel_data[58][6] = 4'b0111; // x=6, y=58
        pixel_data[58][7] = 4'b0111; // x=7, y=58
        pixel_data[58][8] = 4'b0111; // x=8, y=58
        pixel_data[58][9] = 4'b0111; // x=9, y=58
        pixel_data[58][10] = 4'b0111; // x=10, y=58
        pixel_data[58][11] = 4'b0111; // x=11, y=58
        pixel_data[58][12] = 4'b0111; // x=12, y=58
        pixel_data[58][13] = 4'b0111; // x=13, y=58
        pixel_data[58][14] = 4'b0111; // x=14, y=58
        pixel_data[58][15] = 4'b0111; // x=15, y=58
        pixel_data[58][16] = 4'b0111; // x=16, y=58
        pixel_data[58][17] = 4'b0111; // x=17, y=58
        pixel_data[58][18] = 4'b0111; // x=18, y=58
        pixel_data[58][19] = 4'b0111; // x=19, y=58
        pixel_data[58][20] = 4'b0111; // x=20, y=58
        pixel_data[58][21] = 4'b0111; // x=21, y=58
        pixel_data[58][22] = 4'b0111; // x=22, y=58
        pixel_data[58][23] = 4'b0111; // x=23, y=58
        pixel_data[58][24] = 4'b0111; // x=24, y=58
        pixel_data[58][25] = 4'b0111; // x=25, y=58
        pixel_data[58][26] = 4'b0111; // x=26, y=58
        pixel_data[58][27] = 4'b0111; // x=27, y=58
        pixel_data[58][28] = 4'b0111; // x=28, y=58
        pixel_data[58][29] = 4'b0111; // x=29, y=58
        pixel_data[58][30] = 4'b0111; // x=30, y=58
        pixel_data[58][31] = 4'b0111; // x=31, y=58
        pixel_data[58][32] = 4'b0111; // x=32, y=58
        pixel_data[58][33] = 4'b0111; // x=33, y=58
        pixel_data[58][34] = 4'b0111; // x=34, y=58
        pixel_data[58][35] = 4'b0111; // x=35, y=58
        pixel_data[58][36] = 4'b0111; // x=36, y=58
        pixel_data[58][37] = 4'b0111; // x=37, y=58
        pixel_data[58][38] = 4'b0111; // x=38, y=58
        pixel_data[58][39] = 4'b0111; // x=39, y=58
        pixel_data[58][40] = 4'b0111; // x=40, y=58
        pixel_data[58][41] = 4'b0111; // x=41, y=58
        pixel_data[58][42] = 4'b0111; // x=42, y=58
        pixel_data[58][43] = 4'b0111; // x=43, y=58
        pixel_data[58][44] = 4'b0111; // x=44, y=58
        pixel_data[58][45] = 4'b0111; // x=45, y=58
        pixel_data[58][46] = 4'b0111; // x=46, y=58
        pixel_data[58][47] = 4'b0111; // x=47, y=58
        pixel_data[58][48] = 4'b0111; // x=48, y=58
        pixel_data[58][49] = 4'b0111; // x=49, y=58
        pixel_data[58][50] = 4'b0111; // x=50, y=58
        pixel_data[58][51] = 4'b0111; // x=51, y=58
        pixel_data[58][52] = 4'b0111; // x=52, y=58
        pixel_data[58][53] = 4'b0111; // x=53, y=58
        pixel_data[58][54] = 4'b0111; // x=54, y=58
        pixel_data[58][55] = 4'b0111; // x=55, y=58
        pixel_data[58][56] = 4'b0111; // x=56, y=58
        pixel_data[58][57] = 4'b0111; // x=57, y=58
        pixel_data[58][58] = 4'b0111; // x=58, y=58
        pixel_data[58][59] = 4'b0111; // x=59, y=58
        pixel_data[58][60] = 4'b0111; // x=60, y=58
        pixel_data[58][61] = 4'b0111; // x=61, y=58
        pixel_data[58][62] = 4'b0111; // x=62, y=58
        pixel_data[58][63] = 4'b0111; // x=63, y=58
        pixel_data[58][64] = 4'b0111; // x=64, y=58
        pixel_data[58][65] = 4'b0111; // x=65, y=58
        pixel_data[58][66] = 4'b0111; // x=66, y=58
        pixel_data[58][67] = 4'b0111; // x=67, y=58
        pixel_data[58][68] = 4'b0111; // x=68, y=58
        pixel_data[58][69] = 4'b0111; // x=69, y=58
        pixel_data[58][70] = 4'b0111; // x=70, y=58
        pixel_data[58][71] = 4'b0111; // x=71, y=58
        pixel_data[58][72] = 4'b0111; // x=72, y=58
        pixel_data[58][73] = 4'b0111; // x=73, y=58
        pixel_data[58][74] = 4'b0111; // x=74, y=58
        pixel_data[58][75] = 4'b0111; // x=75, y=58
        pixel_data[58][76] = 4'b0111; // x=76, y=58
        pixel_data[58][77] = 4'b0111; // x=77, y=58
        pixel_data[58][78] = 4'b0111; // x=78, y=58
        pixel_data[58][79] = 4'b0111; // x=79, y=58
        pixel_data[58][80] = 4'b0111; // x=80, y=58
        pixel_data[58][81] = 4'b0111; // x=81, y=58
        pixel_data[58][82] = 4'b0111; // x=82, y=58
        pixel_data[58][83] = 4'b0111; // x=83, y=58
        pixel_data[58][84] = 4'b0111; // x=84, y=58
        pixel_data[58][85] = 4'b0111; // x=85, y=58
        pixel_data[58][86] = 4'b0111; // x=86, y=58
        pixel_data[58][87] = 4'b0111; // x=87, y=58
        pixel_data[58][88] = 4'b0111; // x=88, y=58
        pixel_data[58][89] = 4'b0111; // x=89, y=58
        pixel_data[58][90] = 4'b0111; // x=90, y=58
        pixel_data[58][91] = 4'b0111; // x=91, y=58
        pixel_data[58][92] = 4'b0111; // x=92, y=58
        pixel_data[58][93] = 4'b0111; // x=93, y=58
        pixel_data[58][94] = 4'b0111; // x=94, y=58
        pixel_data[58][95] = 4'b0111; // x=95, y=58
        pixel_data[58][96] = 4'b0111; // x=96, y=58
        pixel_data[58][97] = 4'b0111; // x=97, y=58
        pixel_data[58][98] = 4'b0111; // x=98, y=58
        pixel_data[58][99] = 4'b0111; // x=99, y=58
        pixel_data[58][100] = 4'b0111; // x=100, y=58
        pixel_data[58][101] = 4'b0111; // x=101, y=58
        pixel_data[58][102] = 4'b0111; // x=102, y=58
        pixel_data[58][103] = 4'b0111; // x=103, y=58
        pixel_data[58][104] = 4'b0111; // x=104, y=58
        pixel_data[58][105] = 4'b0111; // x=105, y=58
        pixel_data[58][106] = 4'b0111; // x=106, y=58
        pixel_data[58][107] = 4'b0111; // x=107, y=58
        pixel_data[58][108] = 4'b0111; // x=108, y=58
        pixel_data[58][109] = 4'b0111; // x=109, y=58
        pixel_data[58][110] = 4'b0111; // x=110, y=58
        pixel_data[58][111] = 4'b0111; // x=111, y=58
        pixel_data[58][112] = 4'b0111; // x=112, y=58
        pixel_data[58][113] = 4'b0111; // x=113, y=58
        pixel_data[58][114] = 4'b0111; // x=114, y=58
        pixel_data[58][115] = 4'b0111; // x=115, y=58
        pixel_data[58][116] = 4'b0111; // x=116, y=58
        pixel_data[58][117] = 4'b0111; // x=117, y=58
        pixel_data[58][118] = 4'b0111; // x=118, y=58
        pixel_data[58][119] = 4'b0111; // x=119, y=58
        pixel_data[58][120] = 4'b0111; // x=120, y=58
        pixel_data[58][121] = 4'b0111; // x=121, y=58
        pixel_data[58][122] = 4'b0111; // x=122, y=58
        pixel_data[58][123] = 4'b0111; // x=123, y=58
        pixel_data[58][124] = 4'b0111; // x=124, y=58
        pixel_data[58][125] = 4'b0111; // x=125, y=58
        pixel_data[58][126] = 4'b0111; // x=126, y=58
        pixel_data[58][127] = 4'b0111; // x=127, y=58
        pixel_data[58][128] = 4'b0111; // x=128, y=58
        pixel_data[58][129] = 4'b0111; // x=129, y=58
        pixel_data[58][130] = 4'b0111; // x=130, y=58
        pixel_data[58][131] = 4'b0111; // x=131, y=58
        pixel_data[58][132] = 4'b0111; // x=132, y=58
        pixel_data[58][133] = 4'b0111; // x=133, y=58
        pixel_data[58][134] = 4'b0111; // x=134, y=58
        pixel_data[58][135] = 4'b0111; // x=135, y=58
        pixel_data[58][136] = 4'b0111; // x=136, y=58
        pixel_data[58][137] = 4'b0111; // x=137, y=58
        pixel_data[58][138] = 4'b0111; // x=138, y=58
        pixel_data[58][139] = 4'b0111; // x=139, y=58
        pixel_data[58][140] = 4'b0111; // x=140, y=58
        pixel_data[58][141] = 4'b0111; // x=141, y=58
        pixel_data[58][142] = 4'b0111; // x=142, y=58
        pixel_data[58][143] = 4'b0111; // x=143, y=58
        pixel_data[58][144] = 4'b0111; // x=144, y=58
        pixel_data[58][145] = 4'b0111; // x=145, y=58
        pixel_data[58][146] = 4'b0111; // x=146, y=58
        pixel_data[58][147] = 4'b0111; // x=147, y=58
        pixel_data[58][148] = 4'b0111; // x=148, y=58
        pixel_data[58][149] = 4'b0111; // x=149, y=58
        pixel_data[58][150] = 4'b0111; // x=150, y=58
        pixel_data[58][151] = 4'b0111; // x=151, y=58
        pixel_data[58][152] = 4'b0111; // x=152, y=58
        pixel_data[58][153] = 4'b0111; // x=153, y=58
        pixel_data[58][154] = 4'b0111; // x=154, y=58
        pixel_data[58][155] = 4'b0111; // x=155, y=58
        pixel_data[58][156] = 4'b0111; // x=156, y=58
        pixel_data[58][157] = 4'b0111; // x=157, y=58
        pixel_data[58][158] = 4'b0111; // x=158, y=58
        pixel_data[58][159] = 4'b0111; // x=159, y=58
        pixel_data[58][160] = 4'b0111; // x=160, y=58
        pixel_data[58][161] = 4'b0111; // x=161, y=58
        pixel_data[58][162] = 4'b0111; // x=162, y=58
        pixel_data[58][163] = 4'b0111; // x=163, y=58
        pixel_data[58][164] = 4'b0111; // x=164, y=58
        pixel_data[58][165] = 4'b0111; // x=165, y=58
        pixel_data[58][166] = 4'b0111; // x=166, y=58
        pixel_data[58][167] = 4'b0111; // x=167, y=58
        pixel_data[58][168] = 4'b0111; // x=168, y=58
        pixel_data[58][169] = 4'b0111; // x=169, y=58
        pixel_data[58][170] = 4'b0111; // x=170, y=58
        pixel_data[58][171] = 4'b0111; // x=171, y=58
        pixel_data[58][172] = 4'b0111; // x=172, y=58
        pixel_data[58][173] = 4'b0111; // x=173, y=58
        pixel_data[58][174] = 4'b0111; // x=174, y=58
        pixel_data[58][175] = 4'b0111; // x=175, y=58
        pixel_data[58][176] = 4'b0111; // x=176, y=58
        pixel_data[58][177] = 4'b0111; // x=177, y=58
        pixel_data[58][178] = 4'b0111; // x=178, y=58
        pixel_data[58][179] = 4'b0111; // x=179, y=58
        pixel_data[59][0] = 4'b0111; // x=0, y=59
        pixel_data[59][1] = 4'b0111; // x=1, y=59
        pixel_data[59][2] = 4'b0111; // x=2, y=59
        pixel_data[59][3] = 4'b0111; // x=3, y=59
        pixel_data[59][4] = 4'b0111; // x=4, y=59
        pixel_data[59][5] = 4'b0111; // x=5, y=59
        pixel_data[59][6] = 4'b0111; // x=6, y=59
        pixel_data[59][7] = 4'b0111; // x=7, y=59
        pixel_data[59][8] = 4'b0111; // x=8, y=59
        pixel_data[59][9] = 4'b0111; // x=9, y=59
        pixel_data[59][10] = 4'b0111; // x=10, y=59
        pixel_data[59][11] = 4'b0111; // x=11, y=59
        pixel_data[59][12] = 4'b0111; // x=12, y=59
        pixel_data[59][13] = 4'b0111; // x=13, y=59
        pixel_data[59][14] = 4'b0111; // x=14, y=59
        pixel_data[59][15] = 4'b0111; // x=15, y=59
        pixel_data[59][16] = 4'b0111; // x=16, y=59
        pixel_data[59][17] = 4'b0111; // x=17, y=59
        pixel_data[59][18] = 4'b0111; // x=18, y=59
        pixel_data[59][19] = 4'b0111; // x=19, y=59
        pixel_data[59][20] = 4'b0111; // x=20, y=59
        pixel_data[59][21] = 4'b0111; // x=21, y=59
        pixel_data[59][22] = 4'b0111; // x=22, y=59
        pixel_data[59][23] = 4'b0111; // x=23, y=59
        pixel_data[59][24] = 4'b0111; // x=24, y=59
        pixel_data[59][25] = 4'b0111; // x=25, y=59
        pixel_data[59][26] = 4'b0111; // x=26, y=59
        pixel_data[59][27] = 4'b0111; // x=27, y=59
        pixel_data[59][28] = 4'b0111; // x=28, y=59
        pixel_data[59][29] = 4'b0111; // x=29, y=59
        pixel_data[59][30] = 4'b0111; // x=30, y=59
        pixel_data[59][31] = 4'b0111; // x=31, y=59
        pixel_data[59][32] = 4'b0111; // x=32, y=59
        pixel_data[59][33] = 4'b0111; // x=33, y=59
        pixel_data[59][34] = 4'b0111; // x=34, y=59
        pixel_data[59][35] = 4'b0111; // x=35, y=59
        pixel_data[59][36] = 4'b0111; // x=36, y=59
        pixel_data[59][37] = 4'b0111; // x=37, y=59
        pixel_data[59][38] = 4'b0111; // x=38, y=59
        pixel_data[59][39] = 4'b0111; // x=39, y=59
        pixel_data[59][40] = 4'b0111; // x=40, y=59
        pixel_data[59][41] = 4'b0111; // x=41, y=59
        pixel_data[59][42] = 4'b0111; // x=42, y=59
        pixel_data[59][43] = 4'b0111; // x=43, y=59
        pixel_data[59][44] = 4'b0111; // x=44, y=59
        pixel_data[59][45] = 4'b0111; // x=45, y=59
        pixel_data[59][46] = 4'b0111; // x=46, y=59
        pixel_data[59][47] = 4'b0111; // x=47, y=59
        pixel_data[59][48] = 4'b0111; // x=48, y=59
        pixel_data[59][49] = 4'b0111; // x=49, y=59
        pixel_data[59][50] = 4'b0111; // x=50, y=59
        pixel_data[59][51] = 4'b0111; // x=51, y=59
        pixel_data[59][52] = 4'b0111; // x=52, y=59
        pixel_data[59][53] = 4'b0111; // x=53, y=59
        pixel_data[59][54] = 4'b0111; // x=54, y=59
        pixel_data[59][55] = 4'b0111; // x=55, y=59
        pixel_data[59][56] = 4'b0111; // x=56, y=59
        pixel_data[59][57] = 4'b0111; // x=57, y=59
        pixel_data[59][58] = 4'b0111; // x=58, y=59
        pixel_data[59][59] = 4'b0111; // x=59, y=59
        pixel_data[59][60] = 4'b0111; // x=60, y=59
        pixel_data[59][61] = 4'b0111; // x=61, y=59
        pixel_data[59][62] = 4'b0111; // x=62, y=59
        pixel_data[59][63] = 4'b0111; // x=63, y=59
        pixel_data[59][64] = 4'b0111; // x=64, y=59
        pixel_data[59][65] = 4'b0111; // x=65, y=59
        pixel_data[59][66] = 4'b0111; // x=66, y=59
        pixel_data[59][67] = 4'b0111; // x=67, y=59
        pixel_data[59][68] = 4'b0111; // x=68, y=59
        pixel_data[59][69] = 4'b0111; // x=69, y=59
        pixel_data[59][70] = 4'b0111; // x=70, y=59
        pixel_data[59][71] = 4'b0111; // x=71, y=59
        pixel_data[59][72] = 4'b0111; // x=72, y=59
        pixel_data[59][73] = 4'b0111; // x=73, y=59
        pixel_data[59][74] = 4'b0111; // x=74, y=59
        pixel_data[59][75] = 4'b0111; // x=75, y=59
        pixel_data[59][76] = 4'b0111; // x=76, y=59
        pixel_data[59][77] = 4'b0111; // x=77, y=59
        pixel_data[59][78] = 4'b0111; // x=78, y=59
        pixel_data[59][79] = 4'b0111; // x=79, y=59
        pixel_data[59][80] = 4'b0111; // x=80, y=59
        pixel_data[59][81] = 4'b0111; // x=81, y=59
        pixel_data[59][82] = 4'b0111; // x=82, y=59
        pixel_data[59][83] = 4'b0111; // x=83, y=59
        pixel_data[59][84] = 4'b0111; // x=84, y=59
        pixel_data[59][85] = 4'b0111; // x=85, y=59
        pixel_data[59][86] = 4'b0111; // x=86, y=59
        pixel_data[59][87] = 4'b0111; // x=87, y=59
        pixel_data[59][88] = 4'b0111; // x=88, y=59
        pixel_data[59][89] = 4'b0111; // x=89, y=59
        pixel_data[59][90] = 4'b0111; // x=90, y=59
        pixel_data[59][91] = 4'b0111; // x=91, y=59
        pixel_data[59][92] = 4'b0111; // x=92, y=59
        pixel_data[59][93] = 4'b0111; // x=93, y=59
        pixel_data[59][94] = 4'b0111; // x=94, y=59
        pixel_data[59][95] = 4'b0111; // x=95, y=59
        pixel_data[59][96] = 4'b0111; // x=96, y=59
        pixel_data[59][97] = 4'b0111; // x=97, y=59
        pixel_data[59][98] = 4'b0111; // x=98, y=59
        pixel_data[59][99] = 4'b0111; // x=99, y=59
        pixel_data[59][100] = 4'b0111; // x=100, y=59
        pixel_data[59][101] = 4'b0111; // x=101, y=59
        pixel_data[59][102] = 4'b0111; // x=102, y=59
        pixel_data[59][103] = 4'b0111; // x=103, y=59
        pixel_data[59][104] = 4'b0111; // x=104, y=59
        pixel_data[59][105] = 4'b0111; // x=105, y=59
        pixel_data[59][106] = 4'b0111; // x=106, y=59
        pixel_data[59][107] = 4'b0111; // x=107, y=59
        pixel_data[59][108] = 4'b0111; // x=108, y=59
        pixel_data[59][109] = 4'b0111; // x=109, y=59
        pixel_data[59][110] = 4'b0111; // x=110, y=59
        pixel_data[59][111] = 4'b0111; // x=111, y=59
        pixel_data[59][112] = 4'b0111; // x=112, y=59
        pixel_data[59][113] = 4'b0111; // x=113, y=59
        pixel_data[59][114] = 4'b0111; // x=114, y=59
        pixel_data[59][115] = 4'b0111; // x=115, y=59
        pixel_data[59][116] = 4'b0111; // x=116, y=59
        pixel_data[59][117] = 4'b0111; // x=117, y=59
        pixel_data[59][118] = 4'b0111; // x=118, y=59
        pixel_data[59][119] = 4'b0111; // x=119, y=59
        pixel_data[59][120] = 4'b0111; // x=120, y=59
        pixel_data[59][121] = 4'b0111; // x=121, y=59
        pixel_data[59][122] = 4'b0111; // x=122, y=59
        pixel_data[59][123] = 4'b0111; // x=123, y=59
        pixel_data[59][124] = 4'b0111; // x=124, y=59
        pixel_data[59][125] = 4'b0111; // x=125, y=59
        pixel_data[59][126] = 4'b0111; // x=126, y=59
        pixel_data[59][127] = 4'b0111; // x=127, y=59
        pixel_data[59][128] = 4'b0111; // x=128, y=59
        pixel_data[59][129] = 4'b0111; // x=129, y=59
        pixel_data[59][130] = 4'b0111; // x=130, y=59
        pixel_data[59][131] = 4'b0111; // x=131, y=59
        pixel_data[59][132] = 4'b0111; // x=132, y=59
        pixel_data[59][133] = 4'b0111; // x=133, y=59
        pixel_data[59][134] = 4'b0111; // x=134, y=59
        pixel_data[59][135] = 4'b0111; // x=135, y=59
        pixel_data[59][136] = 4'b0111; // x=136, y=59
        pixel_data[59][137] = 4'b0111; // x=137, y=59
        pixel_data[59][138] = 4'b0111; // x=138, y=59
        pixel_data[59][139] = 4'b0111; // x=139, y=59
        pixel_data[59][140] = 4'b0111; // x=140, y=59
        pixel_data[59][141] = 4'b0111; // x=141, y=59
        pixel_data[59][142] = 4'b0111; // x=142, y=59
        pixel_data[59][143] = 4'b0111; // x=143, y=59
        pixel_data[59][144] = 4'b0111; // x=144, y=59
        pixel_data[59][145] = 4'b0111; // x=145, y=59
        pixel_data[59][146] = 4'b0111; // x=146, y=59
        pixel_data[59][147] = 4'b0111; // x=147, y=59
        pixel_data[59][148] = 4'b0111; // x=148, y=59
        pixel_data[59][149] = 4'b0111; // x=149, y=59
        pixel_data[59][150] = 4'b0111; // x=150, y=59
        pixel_data[59][151] = 4'b0111; // x=151, y=59
        pixel_data[59][152] = 4'b0111; // x=152, y=59
        pixel_data[59][153] = 4'b0111; // x=153, y=59
        pixel_data[59][154] = 4'b0111; // x=154, y=59
        pixel_data[59][155] = 4'b0111; // x=155, y=59
        pixel_data[59][156] = 4'b0111; // x=156, y=59
        pixel_data[59][157] = 4'b0111; // x=157, y=59
        pixel_data[59][158] = 4'b0111; // x=158, y=59
        pixel_data[59][159] = 4'b0111; // x=159, y=59
        pixel_data[59][160] = 4'b0111; // x=160, y=59
        pixel_data[59][161] = 4'b0111; // x=161, y=59
        pixel_data[59][162] = 4'b0111; // x=162, y=59
        pixel_data[59][163] = 4'b0111; // x=163, y=59
        pixel_data[59][164] = 4'b0111; // x=164, y=59
        pixel_data[59][165] = 4'b0111; // x=165, y=59
        pixel_data[59][166] = 4'b0111; // x=166, y=59
        pixel_data[59][167] = 4'b0111; // x=167, y=59
        pixel_data[59][168] = 4'b0111; // x=168, y=59
        pixel_data[59][169] = 4'b0111; // x=169, y=59
        pixel_data[59][170] = 4'b0111; // x=170, y=59
        pixel_data[59][171] = 4'b0111; // x=171, y=59
        pixel_data[59][172] = 4'b0111; // x=172, y=59
        pixel_data[59][173] = 4'b0111; // x=173, y=59
        pixel_data[59][174] = 4'b0111; // x=174, y=59
        pixel_data[59][175] = 4'b0111; // x=175, y=59
        pixel_data[59][176] = 4'b0111; // x=176, y=59
        pixel_data[59][177] = 4'b0111; // x=177, y=59
        pixel_data[59][178] = 4'b0111; // x=178, y=59
        pixel_data[59][179] = 4'b0111; // x=179, y=59
    end
endmodule

