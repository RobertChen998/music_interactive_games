module color_palette7(output reg [23:0] color_map [0:15]);
    initial begin
        color_map[0] = 24'hc8c8c8;
        color_map[1] = 24'h000000;
        color_map[2] = 24'hfafafa;
        color_map[3] = 24'h555555;
        color_map[4] = 24'he4e4e4;
        color_map[5] = 24'h909090;
        color_map[6] = 24'h313131;
        color_map[7] = 24'hbdbdbd;
        color_map[8] = 24'h0d0d0d;
        color_map[9] = 24'h616161;
        color_map[10] = 24'hfefefe;
        color_map[11] = 24'h040404;
        color_map[12] = 24'h787878;
        color_map[13] = 24'haaaaaa;
        color_map[14] = 24'h1b1b1b;
        color_map[15] = 24'h454545;
    end
endmodule

module image_data7(output reg [3:0] pixel_data [0:59][0:59]);
    initial begin
        pixel_data[0][0] = 4'b0001; // x=0, y=0
        pixel_data[0][1] = 4'b0001; // x=1, y=0
        pixel_data[0][2] = 4'b0001; // x=2, y=0
        pixel_data[0][3] = 4'b0001; // x=3, y=0
        pixel_data[0][4] = 4'b0001; // x=4, y=0
        pixel_data[0][5] = 4'b0001; // x=5, y=0
        pixel_data[0][6] = 4'b0001; // x=6, y=0
        pixel_data[0][7] = 4'b0001; // x=7, y=0
        pixel_data[0][8] = 4'b0001; // x=8, y=0
        pixel_data[0][9] = 4'b0001; // x=9, y=0
        pixel_data[0][10] = 4'b0001; // x=10, y=0
        pixel_data[0][11] = 4'b0001; // x=11, y=0
        pixel_data[0][12] = 4'b0001; // x=12, y=0
        pixel_data[0][13] = 4'b0001; // x=13, y=0
        pixel_data[0][14] = 4'b0001; // x=14, y=0
        pixel_data[0][15] = 4'b0001; // x=15, y=0
        pixel_data[0][16] = 4'b0001; // x=16, y=0
        pixel_data[0][17] = 4'b0001; // x=17, y=0
        pixel_data[0][18] = 4'b0001; // x=18, y=0
        pixel_data[0][19] = 4'b0001; // x=19, y=0
        pixel_data[0][20] = 4'b0001; // x=20, y=0
        pixel_data[0][21] = 4'b0001; // x=21, y=0
        pixel_data[0][22] = 4'b0001; // x=22, y=0
        pixel_data[0][23] = 4'b0001; // x=23, y=0
        pixel_data[0][24] = 4'b0001; // x=24, y=0
        pixel_data[0][25] = 4'b0001; // x=25, y=0
        pixel_data[0][26] = 4'b0001; // x=26, y=0
        pixel_data[0][27] = 4'b0001; // x=27, y=0
        pixel_data[0][28] = 4'b0001; // x=28, y=0
        pixel_data[0][29] = 4'b0001; // x=29, y=0
        pixel_data[0][30] = 4'b0001; // x=30, y=0
        pixel_data[0][31] = 4'b0001; // x=31, y=0
        pixel_data[0][32] = 4'b0001; // x=32, y=0
        pixel_data[0][33] = 4'b0001; // x=33, y=0
        pixel_data[0][34] = 4'b0001; // x=34, y=0
        pixel_data[0][35] = 4'b0001; // x=35, y=0
        pixel_data[0][36] = 4'b0001; // x=36, y=0
        pixel_data[0][37] = 4'b0001; // x=37, y=0
        pixel_data[0][38] = 4'b0001; // x=38, y=0
        pixel_data[0][39] = 4'b0001; // x=39, y=0
        pixel_data[0][40] = 4'b0001; // x=40, y=0
        pixel_data[0][41] = 4'b0001; // x=41, y=0
        pixel_data[0][42] = 4'b0001; // x=42, y=0
        pixel_data[0][43] = 4'b0001; // x=43, y=0
        pixel_data[0][44] = 4'b0001; // x=44, y=0
        pixel_data[0][45] = 4'b0001; // x=45, y=0
        pixel_data[0][46] = 4'b0001; // x=46, y=0
        pixel_data[0][47] = 4'b0001; // x=47, y=0
        pixel_data[0][48] = 4'b0001; // x=48, y=0
        pixel_data[0][49] = 4'b0001; // x=49, y=0
        pixel_data[0][50] = 4'b0001; // x=50, y=0
        pixel_data[0][51] = 4'b0001; // x=51, y=0
        pixel_data[0][52] = 4'b0001; // x=52, y=0
        pixel_data[0][53] = 4'b0001; // x=53, y=0
        pixel_data[0][54] = 4'b0001; // x=54, y=0
        pixel_data[0][55] = 4'b0001; // x=55, y=0
        pixel_data[0][56] = 4'b0001; // x=56, y=0
        pixel_data[0][57] = 4'b0001; // x=57, y=0
        pixel_data[0][58] = 4'b0001; // x=58, y=0
        pixel_data[0][59] = 4'b0001; // x=59, y=0
        pixel_data[1][0] = 4'b0001; // x=0, y=1
        pixel_data[1][1] = 4'b0001; // x=1, y=1
        pixel_data[1][2] = 4'b0001; // x=2, y=1
        pixel_data[1][3] = 4'b0001; // x=3, y=1
        pixel_data[1][4] = 4'b0001; // x=4, y=1
        pixel_data[1][5] = 4'b0001; // x=5, y=1
        pixel_data[1][6] = 4'b0001; // x=6, y=1
        pixel_data[1][7] = 4'b0001; // x=7, y=1
        pixel_data[1][8] = 4'b0001; // x=8, y=1
        pixel_data[1][9] = 4'b0001; // x=9, y=1
        pixel_data[1][10] = 4'b0001; // x=10, y=1
        pixel_data[1][11] = 4'b0001; // x=11, y=1
        pixel_data[1][12] = 4'b0001; // x=12, y=1
        pixel_data[1][13] = 4'b0001; // x=13, y=1
        pixel_data[1][14] = 4'b0001; // x=14, y=1
        pixel_data[1][15] = 4'b0001; // x=15, y=1
        pixel_data[1][16] = 4'b0001; // x=16, y=1
        pixel_data[1][17] = 4'b0001; // x=17, y=1
        pixel_data[1][18] = 4'b0001; // x=18, y=1
        pixel_data[1][19] = 4'b0001; // x=19, y=1
        pixel_data[1][20] = 4'b0001; // x=20, y=1
        pixel_data[1][21] = 4'b0001; // x=21, y=1
        pixel_data[1][22] = 4'b0001; // x=22, y=1
        pixel_data[1][23] = 4'b0001; // x=23, y=1
        pixel_data[1][24] = 4'b0001; // x=24, y=1
        pixel_data[1][25] = 4'b0001; // x=25, y=1
        pixel_data[1][26] = 4'b0001; // x=26, y=1
        pixel_data[1][27] = 4'b0001; // x=27, y=1
        pixel_data[1][28] = 4'b0001; // x=28, y=1
        pixel_data[1][29] = 4'b0001; // x=29, y=1
        pixel_data[1][30] = 4'b0001; // x=30, y=1
        pixel_data[1][31] = 4'b0001; // x=31, y=1
        pixel_data[1][32] = 4'b0001; // x=32, y=1
        pixel_data[1][33] = 4'b0001; // x=33, y=1
        pixel_data[1][34] = 4'b0001; // x=34, y=1
        pixel_data[1][35] = 4'b0001; // x=35, y=1
        pixel_data[1][36] = 4'b0001; // x=36, y=1
        pixel_data[1][37] = 4'b0001; // x=37, y=1
        pixel_data[1][38] = 4'b0001; // x=38, y=1
        pixel_data[1][39] = 4'b0001; // x=39, y=1
        pixel_data[1][40] = 4'b0001; // x=40, y=1
        pixel_data[1][41] = 4'b0001; // x=41, y=1
        pixel_data[1][42] = 4'b0001; // x=42, y=1
        pixel_data[1][43] = 4'b0001; // x=43, y=1
        pixel_data[1][44] = 4'b0001; // x=44, y=1
        pixel_data[1][45] = 4'b0001; // x=45, y=1
        pixel_data[1][46] = 4'b0001; // x=46, y=1
        pixel_data[1][47] = 4'b0001; // x=47, y=1
        pixel_data[1][48] = 4'b0001; // x=48, y=1
        pixel_data[1][49] = 4'b0001; // x=49, y=1
        pixel_data[1][50] = 4'b0001; // x=50, y=1
        pixel_data[1][51] = 4'b0001; // x=51, y=1
        pixel_data[1][52] = 4'b0001; // x=52, y=1
        pixel_data[1][53] = 4'b0001; // x=53, y=1
        pixel_data[1][54] = 4'b0001; // x=54, y=1
        pixel_data[1][55] = 4'b0001; // x=55, y=1
        pixel_data[1][56] = 4'b0001; // x=56, y=1
        pixel_data[1][57] = 4'b0001; // x=57, y=1
        pixel_data[1][58] = 4'b0001; // x=58, y=1
        pixel_data[1][59] = 4'b0001; // x=59, y=1
        pixel_data[2][0] = 4'b0001; // x=0, y=2
        pixel_data[2][1] = 4'b0001; // x=1, y=2
        pixel_data[2][2] = 4'b0001; // x=2, y=2
        pixel_data[2][3] = 4'b0001; // x=3, y=2
        pixel_data[2][4] = 4'b0001; // x=4, y=2
        pixel_data[2][5] = 4'b0001; // x=5, y=2
        pixel_data[2][6] = 4'b0001; // x=6, y=2
        pixel_data[2][7] = 4'b0001; // x=7, y=2
        pixel_data[2][8] = 4'b0001; // x=8, y=2
        pixel_data[2][9] = 4'b0001; // x=9, y=2
        pixel_data[2][10] = 4'b0001; // x=10, y=2
        pixel_data[2][11] = 4'b0001; // x=11, y=2
        pixel_data[2][12] = 4'b0001; // x=12, y=2
        pixel_data[2][13] = 4'b0001; // x=13, y=2
        pixel_data[2][14] = 4'b0001; // x=14, y=2
        pixel_data[2][15] = 4'b0001; // x=15, y=2
        pixel_data[2][16] = 4'b0001; // x=16, y=2
        pixel_data[2][17] = 4'b0001; // x=17, y=2
        pixel_data[2][18] = 4'b0001; // x=18, y=2
        pixel_data[2][19] = 4'b0001; // x=19, y=2
        pixel_data[2][20] = 4'b0001; // x=20, y=2
        pixel_data[2][21] = 4'b0001; // x=21, y=2
        pixel_data[2][22] = 4'b0001; // x=22, y=2
        pixel_data[2][23] = 4'b0001; // x=23, y=2
        pixel_data[2][24] = 4'b0001; // x=24, y=2
        pixel_data[2][25] = 4'b0001; // x=25, y=2
        pixel_data[2][26] = 4'b0001; // x=26, y=2
        pixel_data[2][27] = 4'b0001; // x=27, y=2
        pixel_data[2][28] = 4'b0001; // x=28, y=2
        pixel_data[2][29] = 4'b0001; // x=29, y=2
        pixel_data[2][30] = 4'b0001; // x=30, y=2
        pixel_data[2][31] = 4'b0001; // x=31, y=2
        pixel_data[2][32] = 4'b0001; // x=32, y=2
        pixel_data[2][33] = 4'b0001; // x=33, y=2
        pixel_data[2][34] = 4'b0001; // x=34, y=2
        pixel_data[2][35] = 4'b0001; // x=35, y=2
        pixel_data[2][36] = 4'b0001; // x=36, y=2
        pixel_data[2][37] = 4'b0001; // x=37, y=2
        pixel_data[2][38] = 4'b0001; // x=38, y=2
        pixel_data[2][39] = 4'b0001; // x=39, y=2
        pixel_data[2][40] = 4'b0001; // x=40, y=2
        pixel_data[2][41] = 4'b0001; // x=41, y=2
        pixel_data[2][42] = 4'b0001; // x=42, y=2
        pixel_data[2][43] = 4'b0001; // x=43, y=2
        pixel_data[2][44] = 4'b0001; // x=44, y=2
        pixel_data[2][45] = 4'b0001; // x=45, y=2
        pixel_data[2][46] = 4'b0001; // x=46, y=2
        pixel_data[2][47] = 4'b0001; // x=47, y=2
        pixel_data[2][48] = 4'b0001; // x=48, y=2
        pixel_data[2][49] = 4'b0001; // x=49, y=2
        pixel_data[2][50] = 4'b0001; // x=50, y=2
        pixel_data[2][51] = 4'b0001; // x=51, y=2
        pixel_data[2][52] = 4'b0001; // x=52, y=2
        pixel_data[2][53] = 4'b0001; // x=53, y=2
        pixel_data[2][54] = 4'b0001; // x=54, y=2
        pixel_data[2][55] = 4'b0001; // x=55, y=2
        pixel_data[2][56] = 4'b0001; // x=56, y=2
        pixel_data[2][57] = 4'b0001; // x=57, y=2
        pixel_data[2][58] = 4'b0001; // x=58, y=2
        pixel_data[2][59] = 4'b0001; // x=59, y=2
        pixel_data[3][0] = 4'b0001; // x=0, y=3
        pixel_data[3][1] = 4'b0001; // x=1, y=3
        pixel_data[3][2] = 4'b0001; // x=2, y=3
        pixel_data[3][3] = 4'b0001; // x=3, y=3
        pixel_data[3][4] = 4'b0001; // x=4, y=3
        pixel_data[3][5] = 4'b0001; // x=5, y=3
        pixel_data[3][6] = 4'b0001; // x=6, y=3
        pixel_data[3][7] = 4'b0001; // x=7, y=3
        pixel_data[3][8] = 4'b0001; // x=8, y=3
        pixel_data[3][9] = 4'b0001; // x=9, y=3
        pixel_data[3][10] = 4'b0001; // x=10, y=3
        pixel_data[3][11] = 4'b0001; // x=11, y=3
        pixel_data[3][12] = 4'b0001; // x=12, y=3
        pixel_data[3][13] = 4'b0001; // x=13, y=3
        pixel_data[3][14] = 4'b0001; // x=14, y=3
        pixel_data[3][15] = 4'b0001; // x=15, y=3
        pixel_data[3][16] = 4'b0001; // x=16, y=3
        pixel_data[3][17] = 4'b0001; // x=17, y=3
        pixel_data[3][18] = 4'b0001; // x=18, y=3
        pixel_data[3][19] = 4'b0001; // x=19, y=3
        pixel_data[3][20] = 4'b0001; // x=20, y=3
        pixel_data[3][21] = 4'b0001; // x=21, y=3
        pixel_data[3][22] = 4'b0001; // x=22, y=3
        pixel_data[3][23] = 4'b0001; // x=23, y=3
        pixel_data[3][24] = 4'b0001; // x=24, y=3
        pixel_data[3][25] = 4'b0001; // x=25, y=3
        pixel_data[3][26] = 4'b0001; // x=26, y=3
        pixel_data[3][27] = 4'b0001; // x=27, y=3
        pixel_data[3][28] = 4'b0001; // x=28, y=3
        pixel_data[3][29] = 4'b0001; // x=29, y=3
        pixel_data[3][30] = 4'b0001; // x=30, y=3
        pixel_data[3][31] = 4'b0001; // x=31, y=3
        pixel_data[3][32] = 4'b0001; // x=32, y=3
        pixel_data[3][33] = 4'b0001; // x=33, y=3
        pixel_data[3][34] = 4'b0001; // x=34, y=3
        pixel_data[3][35] = 4'b0001; // x=35, y=3
        pixel_data[3][36] = 4'b0001; // x=36, y=3
        pixel_data[3][37] = 4'b0001; // x=37, y=3
        pixel_data[3][38] = 4'b0001; // x=38, y=3
        pixel_data[3][39] = 4'b0001; // x=39, y=3
        pixel_data[3][40] = 4'b0001; // x=40, y=3
        pixel_data[3][41] = 4'b0001; // x=41, y=3
        pixel_data[3][42] = 4'b0001; // x=42, y=3
        pixel_data[3][43] = 4'b0001; // x=43, y=3
        pixel_data[3][44] = 4'b0001; // x=44, y=3
        pixel_data[3][45] = 4'b0001; // x=45, y=3
        pixel_data[3][46] = 4'b0001; // x=46, y=3
        pixel_data[3][47] = 4'b0001; // x=47, y=3
        pixel_data[3][48] = 4'b0001; // x=48, y=3
        pixel_data[3][49] = 4'b0001; // x=49, y=3
        pixel_data[3][50] = 4'b0001; // x=50, y=3
        pixel_data[3][51] = 4'b0001; // x=51, y=3
        pixel_data[3][52] = 4'b0001; // x=52, y=3
        pixel_data[3][53] = 4'b0001; // x=53, y=3
        pixel_data[3][54] = 4'b0001; // x=54, y=3
        pixel_data[3][55] = 4'b0001; // x=55, y=3
        pixel_data[3][56] = 4'b0001; // x=56, y=3
        pixel_data[3][57] = 4'b0001; // x=57, y=3
        pixel_data[3][58] = 4'b0001; // x=58, y=3
        pixel_data[3][59] = 4'b0001; // x=59, y=3
        pixel_data[4][0] = 4'b0001; // x=0, y=4
        pixel_data[4][1] = 4'b0001; // x=1, y=4
        pixel_data[4][2] = 4'b0001; // x=2, y=4
        pixel_data[4][3] = 4'b0001; // x=3, y=4
        pixel_data[4][4] = 4'b0001; // x=4, y=4
        pixel_data[4][5] = 4'b0001; // x=5, y=4
        pixel_data[4][6] = 4'b0001; // x=6, y=4
        pixel_data[4][7] = 4'b0001; // x=7, y=4
        pixel_data[4][8] = 4'b0001; // x=8, y=4
        pixel_data[4][9] = 4'b0001; // x=9, y=4
        pixel_data[4][10] = 4'b0001; // x=10, y=4
        pixel_data[4][11] = 4'b0001; // x=11, y=4
        pixel_data[4][12] = 4'b0001; // x=12, y=4
        pixel_data[4][13] = 4'b0001; // x=13, y=4
        pixel_data[4][14] = 4'b0001; // x=14, y=4
        pixel_data[4][15] = 4'b0001; // x=15, y=4
        pixel_data[4][16] = 4'b0001; // x=16, y=4
        pixel_data[4][17] = 4'b0001; // x=17, y=4
        pixel_data[4][18] = 4'b0001; // x=18, y=4
        pixel_data[4][19] = 4'b0001; // x=19, y=4
        pixel_data[4][20] = 4'b0001; // x=20, y=4
        pixel_data[4][21] = 4'b0001; // x=21, y=4
        pixel_data[4][22] = 4'b0001; // x=22, y=4
        pixel_data[4][23] = 4'b0001; // x=23, y=4
        pixel_data[4][24] = 4'b0001; // x=24, y=4
        pixel_data[4][25] = 4'b0001; // x=25, y=4
        pixel_data[4][26] = 4'b0001; // x=26, y=4
        pixel_data[4][27] = 4'b0001; // x=27, y=4
        pixel_data[4][28] = 4'b0001; // x=28, y=4
        pixel_data[4][29] = 4'b0001; // x=29, y=4
        pixel_data[4][30] = 4'b0001; // x=30, y=4
        pixel_data[4][31] = 4'b0001; // x=31, y=4
        pixel_data[4][32] = 4'b0001; // x=32, y=4
        pixel_data[4][33] = 4'b0001; // x=33, y=4
        pixel_data[4][34] = 4'b0001; // x=34, y=4
        pixel_data[4][35] = 4'b0001; // x=35, y=4
        pixel_data[4][36] = 4'b0001; // x=36, y=4
        pixel_data[4][37] = 4'b0001; // x=37, y=4
        pixel_data[4][38] = 4'b0001; // x=38, y=4
        pixel_data[4][39] = 4'b0001; // x=39, y=4
        pixel_data[4][40] = 4'b0001; // x=40, y=4
        pixel_data[4][41] = 4'b0001; // x=41, y=4
        pixel_data[4][42] = 4'b0001; // x=42, y=4
        pixel_data[4][43] = 4'b0001; // x=43, y=4
        pixel_data[4][44] = 4'b0001; // x=44, y=4
        pixel_data[4][45] = 4'b0001; // x=45, y=4
        pixel_data[4][46] = 4'b0001; // x=46, y=4
        pixel_data[4][47] = 4'b0001; // x=47, y=4
        pixel_data[4][48] = 4'b0001; // x=48, y=4
        pixel_data[4][49] = 4'b0001; // x=49, y=4
        pixel_data[4][50] = 4'b0001; // x=50, y=4
        pixel_data[4][51] = 4'b0001; // x=51, y=4
        pixel_data[4][52] = 4'b0001; // x=52, y=4
        pixel_data[4][53] = 4'b0001; // x=53, y=4
        pixel_data[4][54] = 4'b0001; // x=54, y=4
        pixel_data[4][55] = 4'b0001; // x=55, y=4
        pixel_data[4][56] = 4'b0001; // x=56, y=4
        pixel_data[4][57] = 4'b0001; // x=57, y=4
        pixel_data[4][58] = 4'b0001; // x=58, y=4
        pixel_data[4][59] = 4'b0001; // x=59, y=4
        pixel_data[5][0] = 4'b0001; // x=0, y=5
        pixel_data[5][1] = 4'b0001; // x=1, y=5
        pixel_data[5][2] = 4'b0001; // x=2, y=5
        pixel_data[5][3] = 4'b0001; // x=3, y=5
        pixel_data[5][4] = 4'b0001; // x=4, y=5
        pixel_data[5][5] = 4'b0001; // x=5, y=5
        pixel_data[5][6] = 4'b0001; // x=6, y=5
        pixel_data[5][7] = 4'b0001; // x=7, y=5
        pixel_data[5][8] = 4'b0001; // x=8, y=5
        pixel_data[5][9] = 4'b0001; // x=9, y=5
        pixel_data[5][10] = 4'b0001; // x=10, y=5
        pixel_data[5][11] = 4'b0001; // x=11, y=5
        pixel_data[5][12] = 4'b0001; // x=12, y=5
        pixel_data[5][13] = 4'b0001; // x=13, y=5
        pixel_data[5][14] = 4'b0001; // x=14, y=5
        pixel_data[5][15] = 4'b0001; // x=15, y=5
        pixel_data[5][16] = 4'b0001; // x=16, y=5
        pixel_data[5][17] = 4'b0001; // x=17, y=5
        pixel_data[5][18] = 4'b0001; // x=18, y=5
        pixel_data[5][19] = 4'b0001; // x=19, y=5
        pixel_data[5][20] = 4'b0001; // x=20, y=5
        pixel_data[5][21] = 4'b0001; // x=21, y=5
        pixel_data[5][22] = 4'b0001; // x=22, y=5
        pixel_data[5][23] = 4'b0001; // x=23, y=5
        pixel_data[5][24] = 4'b0001; // x=24, y=5
        pixel_data[5][25] = 4'b0001; // x=25, y=5
        pixel_data[5][26] = 4'b0001; // x=26, y=5
        pixel_data[5][27] = 4'b0001; // x=27, y=5
        pixel_data[5][28] = 4'b0001; // x=28, y=5
        pixel_data[5][29] = 4'b0001; // x=29, y=5
        pixel_data[5][30] = 4'b0001; // x=30, y=5
        pixel_data[5][31] = 4'b0001; // x=31, y=5
        pixel_data[5][32] = 4'b0001; // x=32, y=5
        pixel_data[5][33] = 4'b0001; // x=33, y=5
        pixel_data[5][34] = 4'b0001; // x=34, y=5
        pixel_data[5][35] = 4'b0001; // x=35, y=5
        pixel_data[5][36] = 4'b0001; // x=36, y=5
        pixel_data[5][37] = 4'b0001; // x=37, y=5
        pixel_data[5][38] = 4'b0001; // x=38, y=5
        pixel_data[5][39] = 4'b0001; // x=39, y=5
        pixel_data[5][40] = 4'b0001; // x=40, y=5
        pixel_data[5][41] = 4'b0001; // x=41, y=5
        pixel_data[5][42] = 4'b0001; // x=42, y=5
        pixel_data[5][43] = 4'b0001; // x=43, y=5
        pixel_data[5][44] = 4'b0001; // x=44, y=5
        pixel_data[5][45] = 4'b0001; // x=45, y=5
        pixel_data[5][46] = 4'b0001; // x=46, y=5
        pixel_data[5][47] = 4'b0001; // x=47, y=5
        pixel_data[5][48] = 4'b0001; // x=48, y=5
        pixel_data[5][49] = 4'b0001; // x=49, y=5
        pixel_data[5][50] = 4'b0001; // x=50, y=5
        pixel_data[5][51] = 4'b0001; // x=51, y=5
        pixel_data[5][52] = 4'b0001; // x=52, y=5
        pixel_data[5][53] = 4'b0001; // x=53, y=5
        pixel_data[5][54] = 4'b0001; // x=54, y=5
        pixel_data[5][55] = 4'b0001; // x=55, y=5
        pixel_data[5][56] = 4'b0001; // x=56, y=5
        pixel_data[5][57] = 4'b0001; // x=57, y=5
        pixel_data[5][58] = 4'b0001; // x=58, y=5
        pixel_data[5][59] = 4'b0001; // x=59, y=5
        pixel_data[6][0] = 4'b0001; // x=0, y=6
        pixel_data[6][1] = 4'b0001; // x=1, y=6
        pixel_data[6][2] = 4'b0001; // x=2, y=6
        pixel_data[6][3] = 4'b0001; // x=3, y=6
        pixel_data[6][4] = 4'b0001; // x=4, y=6
        pixel_data[6][5] = 4'b0001; // x=5, y=6
        pixel_data[6][6] = 4'b0001; // x=6, y=6
        pixel_data[6][7] = 4'b0001; // x=7, y=6
        pixel_data[6][8] = 4'b0001; // x=8, y=6
        pixel_data[6][9] = 4'b0001; // x=9, y=6
        pixel_data[6][10] = 4'b0001; // x=10, y=6
        pixel_data[6][11] = 4'b0001; // x=11, y=6
        pixel_data[6][12] = 4'b0001; // x=12, y=6
        pixel_data[6][13] = 4'b0001; // x=13, y=6
        pixel_data[6][14] = 4'b0001; // x=14, y=6
        pixel_data[6][15] = 4'b0001; // x=15, y=6
        pixel_data[6][16] = 4'b0001; // x=16, y=6
        pixel_data[6][17] = 4'b0001; // x=17, y=6
        pixel_data[6][18] = 4'b0001; // x=18, y=6
        pixel_data[6][19] = 4'b0001; // x=19, y=6
        pixel_data[6][20] = 4'b0001; // x=20, y=6
        pixel_data[6][21] = 4'b0001; // x=21, y=6
        pixel_data[6][22] = 4'b0001; // x=22, y=6
        pixel_data[6][23] = 4'b0001; // x=23, y=6
        pixel_data[6][24] = 4'b0001; // x=24, y=6
        pixel_data[6][25] = 4'b0001; // x=25, y=6
        pixel_data[6][26] = 4'b0001; // x=26, y=6
        pixel_data[6][27] = 4'b0001; // x=27, y=6
        pixel_data[6][28] = 4'b0001; // x=28, y=6
        pixel_data[6][29] = 4'b0001; // x=29, y=6
        pixel_data[6][30] = 4'b0001; // x=30, y=6
        pixel_data[6][31] = 4'b0001; // x=31, y=6
        pixel_data[6][32] = 4'b0001; // x=32, y=6
        pixel_data[6][33] = 4'b0001; // x=33, y=6
        pixel_data[6][34] = 4'b0001; // x=34, y=6
        pixel_data[6][35] = 4'b0001; // x=35, y=6
        pixel_data[6][36] = 4'b0001; // x=36, y=6
        pixel_data[6][37] = 4'b0001; // x=37, y=6
        pixel_data[6][38] = 4'b0001; // x=38, y=6
        pixel_data[6][39] = 4'b0001; // x=39, y=6
        pixel_data[6][40] = 4'b0001; // x=40, y=6
        pixel_data[6][41] = 4'b0001; // x=41, y=6
        pixel_data[6][42] = 4'b0001; // x=42, y=6
        pixel_data[6][43] = 4'b0001; // x=43, y=6
        pixel_data[6][44] = 4'b0001; // x=44, y=6
        pixel_data[6][45] = 4'b0001; // x=45, y=6
        pixel_data[6][46] = 4'b0001; // x=46, y=6
        pixel_data[6][47] = 4'b0001; // x=47, y=6
        pixel_data[6][48] = 4'b0001; // x=48, y=6
        pixel_data[6][49] = 4'b0001; // x=49, y=6
        pixel_data[6][50] = 4'b0001; // x=50, y=6
        pixel_data[6][51] = 4'b0001; // x=51, y=6
        pixel_data[6][52] = 4'b0001; // x=52, y=6
        pixel_data[6][53] = 4'b0001; // x=53, y=6
        pixel_data[6][54] = 4'b0001; // x=54, y=6
        pixel_data[6][55] = 4'b0001; // x=55, y=6
        pixel_data[6][56] = 4'b0001; // x=56, y=6
        pixel_data[6][57] = 4'b0001; // x=57, y=6
        pixel_data[6][58] = 4'b0001; // x=58, y=6
        pixel_data[6][59] = 4'b0001; // x=59, y=6
        pixel_data[7][0] = 4'b0001; // x=0, y=7
        pixel_data[7][1] = 4'b0001; // x=1, y=7
        pixel_data[7][2] = 4'b0001; // x=2, y=7
        pixel_data[7][3] = 4'b0001; // x=3, y=7
        pixel_data[7][4] = 4'b0001; // x=4, y=7
        pixel_data[7][5] = 4'b0001; // x=5, y=7
        pixel_data[7][6] = 4'b0001; // x=6, y=7
        pixel_data[7][7] = 4'b0001; // x=7, y=7
        pixel_data[7][8] = 4'b0001; // x=8, y=7
        pixel_data[7][9] = 4'b0001; // x=9, y=7
        pixel_data[7][10] = 4'b0001; // x=10, y=7
        pixel_data[7][11] = 4'b0001; // x=11, y=7
        pixel_data[7][12] = 4'b0001; // x=12, y=7
        pixel_data[7][13] = 4'b0001; // x=13, y=7
        pixel_data[7][14] = 4'b0001; // x=14, y=7
        pixel_data[7][15] = 4'b0001; // x=15, y=7
        pixel_data[7][16] = 4'b0001; // x=16, y=7
        pixel_data[7][17] = 4'b0001; // x=17, y=7
        pixel_data[7][18] = 4'b0001; // x=18, y=7
        pixel_data[7][19] = 4'b0001; // x=19, y=7
        pixel_data[7][20] = 4'b0001; // x=20, y=7
        pixel_data[7][21] = 4'b0001; // x=21, y=7
        pixel_data[7][22] = 4'b0001; // x=22, y=7
        pixel_data[7][23] = 4'b0001; // x=23, y=7
        pixel_data[7][24] = 4'b0001; // x=24, y=7
        pixel_data[7][25] = 4'b0001; // x=25, y=7
        pixel_data[7][26] = 4'b0001; // x=26, y=7
        pixel_data[7][27] = 4'b0001; // x=27, y=7
        pixel_data[7][28] = 4'b0001; // x=28, y=7
        pixel_data[7][29] = 4'b0001; // x=29, y=7
        pixel_data[7][30] = 4'b0001; // x=30, y=7
        pixel_data[7][31] = 4'b0001; // x=31, y=7
        pixel_data[7][32] = 4'b0001; // x=32, y=7
        pixel_data[7][33] = 4'b0001; // x=33, y=7
        pixel_data[7][34] = 4'b0001; // x=34, y=7
        pixel_data[7][35] = 4'b0001; // x=35, y=7
        pixel_data[7][36] = 4'b0001; // x=36, y=7
        pixel_data[7][37] = 4'b0001; // x=37, y=7
        pixel_data[7][38] = 4'b0001; // x=38, y=7
        pixel_data[7][39] = 4'b0001; // x=39, y=7
        pixel_data[7][40] = 4'b0001; // x=40, y=7
        pixel_data[7][41] = 4'b0001; // x=41, y=7
        pixel_data[7][42] = 4'b0001; // x=42, y=7
        pixel_data[7][43] = 4'b0001; // x=43, y=7
        pixel_data[7][44] = 4'b0001; // x=44, y=7
        pixel_data[7][45] = 4'b0001; // x=45, y=7
        pixel_data[7][46] = 4'b0001; // x=46, y=7
        pixel_data[7][47] = 4'b0001; // x=47, y=7
        pixel_data[7][48] = 4'b0001; // x=48, y=7
        pixel_data[7][49] = 4'b0001; // x=49, y=7
        pixel_data[7][50] = 4'b0001; // x=50, y=7
        pixel_data[7][51] = 4'b0001; // x=51, y=7
        pixel_data[7][52] = 4'b0001; // x=52, y=7
        pixel_data[7][53] = 4'b0001; // x=53, y=7
        pixel_data[7][54] = 4'b0001; // x=54, y=7
        pixel_data[7][55] = 4'b0001; // x=55, y=7
        pixel_data[7][56] = 4'b0001; // x=56, y=7
        pixel_data[7][57] = 4'b0001; // x=57, y=7
        pixel_data[7][58] = 4'b0001; // x=58, y=7
        pixel_data[7][59] = 4'b0001; // x=59, y=7
        pixel_data[8][0] = 4'b0001; // x=0, y=8
        pixel_data[8][1] = 4'b0001; // x=1, y=8
        pixel_data[8][2] = 4'b0001; // x=2, y=8
        pixel_data[8][3] = 4'b0001; // x=3, y=8
        pixel_data[8][4] = 4'b0001; // x=4, y=8
        pixel_data[8][5] = 4'b0001; // x=5, y=8
        pixel_data[8][6] = 4'b0001; // x=6, y=8
        pixel_data[8][7] = 4'b0001; // x=7, y=8
        pixel_data[8][8] = 4'b0001; // x=8, y=8
        pixel_data[8][9] = 4'b0001; // x=9, y=8
        pixel_data[8][10] = 4'b0001; // x=10, y=8
        pixel_data[8][11] = 4'b0001; // x=11, y=8
        pixel_data[8][12] = 4'b0001; // x=12, y=8
        pixel_data[8][13] = 4'b0001; // x=13, y=8
        pixel_data[8][14] = 4'b0001; // x=14, y=8
        pixel_data[8][15] = 4'b0001; // x=15, y=8
        pixel_data[8][16] = 4'b0001; // x=16, y=8
        pixel_data[8][17] = 4'b0001; // x=17, y=8
        pixel_data[8][18] = 4'b0001; // x=18, y=8
        pixel_data[8][19] = 4'b0001; // x=19, y=8
        pixel_data[8][20] = 4'b0001; // x=20, y=8
        pixel_data[8][21] = 4'b0001; // x=21, y=8
        pixel_data[8][22] = 4'b0001; // x=22, y=8
        pixel_data[8][23] = 4'b0001; // x=23, y=8
        pixel_data[8][24] = 4'b0001; // x=24, y=8
        pixel_data[8][25] = 4'b0001; // x=25, y=8
        pixel_data[8][26] = 4'b0001; // x=26, y=8
        pixel_data[8][27] = 4'b0001; // x=27, y=8
        pixel_data[8][28] = 4'b0001; // x=28, y=8
        pixel_data[8][29] = 4'b0001; // x=29, y=8
        pixel_data[8][30] = 4'b0001; // x=30, y=8
        pixel_data[8][31] = 4'b0001; // x=31, y=8
        pixel_data[8][32] = 4'b0001; // x=32, y=8
        pixel_data[8][33] = 4'b0001; // x=33, y=8
        pixel_data[8][34] = 4'b0001; // x=34, y=8
        pixel_data[8][35] = 4'b0001; // x=35, y=8
        pixel_data[8][36] = 4'b0001; // x=36, y=8
        pixel_data[8][37] = 4'b0001; // x=37, y=8
        pixel_data[8][38] = 4'b0001; // x=38, y=8
        pixel_data[8][39] = 4'b0001; // x=39, y=8
        pixel_data[8][40] = 4'b0001; // x=40, y=8
        pixel_data[8][41] = 4'b0001; // x=41, y=8
        pixel_data[8][42] = 4'b0001; // x=42, y=8
        pixel_data[8][43] = 4'b0001; // x=43, y=8
        pixel_data[8][44] = 4'b0001; // x=44, y=8
        pixel_data[8][45] = 4'b0001; // x=45, y=8
        pixel_data[8][46] = 4'b0001; // x=46, y=8
        pixel_data[8][47] = 4'b0001; // x=47, y=8
        pixel_data[8][48] = 4'b0001; // x=48, y=8
        pixel_data[8][49] = 4'b0001; // x=49, y=8
        pixel_data[8][50] = 4'b0001; // x=50, y=8
        pixel_data[8][51] = 4'b0001; // x=51, y=8
        pixel_data[8][52] = 4'b0001; // x=52, y=8
        pixel_data[8][53] = 4'b0001; // x=53, y=8
        pixel_data[8][54] = 4'b0001; // x=54, y=8
        pixel_data[8][55] = 4'b0001; // x=55, y=8
        pixel_data[8][56] = 4'b0001; // x=56, y=8
        pixel_data[8][57] = 4'b0001; // x=57, y=8
        pixel_data[8][58] = 4'b0001; // x=58, y=8
        pixel_data[8][59] = 4'b0001; // x=59, y=8
        pixel_data[9][0] = 4'b0001; // x=0, y=9
        pixel_data[9][1] = 4'b0001; // x=1, y=9
        pixel_data[9][2] = 4'b0001; // x=2, y=9
        pixel_data[9][3] = 4'b0001; // x=3, y=9
        pixel_data[9][4] = 4'b0001; // x=4, y=9
        pixel_data[9][5] = 4'b0001; // x=5, y=9
        pixel_data[9][6] = 4'b0001; // x=6, y=9
        pixel_data[9][7] = 4'b0001; // x=7, y=9
        pixel_data[9][8] = 4'b0001; // x=8, y=9
        pixel_data[9][9] = 4'b0001; // x=9, y=9
        pixel_data[9][10] = 4'b0001; // x=10, y=9
        pixel_data[9][11] = 4'b0001; // x=11, y=9
        pixel_data[9][12] = 4'b0001; // x=12, y=9
        pixel_data[9][13] = 4'b0001; // x=13, y=9
        pixel_data[9][14] = 4'b0001; // x=14, y=9
        pixel_data[9][15] = 4'b0001; // x=15, y=9
        pixel_data[9][16] = 4'b0001; // x=16, y=9
        pixel_data[9][17] = 4'b0001; // x=17, y=9
        pixel_data[9][18] = 4'b0001; // x=18, y=9
        pixel_data[9][19] = 4'b0001; // x=19, y=9
        pixel_data[9][20] = 4'b0001; // x=20, y=9
        pixel_data[9][21] = 4'b0001; // x=21, y=9
        pixel_data[9][22] = 4'b0001; // x=22, y=9
        pixel_data[9][23] = 4'b0001; // x=23, y=9
        pixel_data[9][24] = 4'b0001; // x=24, y=9
        pixel_data[9][25] = 4'b0001; // x=25, y=9
        pixel_data[9][26] = 4'b0001; // x=26, y=9
        pixel_data[9][27] = 4'b0001; // x=27, y=9
        pixel_data[9][28] = 4'b0001; // x=28, y=9
        pixel_data[9][29] = 4'b0001; // x=29, y=9
        pixel_data[9][30] = 4'b0001; // x=30, y=9
        pixel_data[9][31] = 4'b0001; // x=31, y=9
        pixel_data[9][32] = 4'b0001; // x=32, y=9
        pixel_data[9][33] = 4'b0001; // x=33, y=9
        pixel_data[9][34] = 4'b0001; // x=34, y=9
        pixel_data[9][35] = 4'b0001; // x=35, y=9
        pixel_data[9][36] = 4'b0001; // x=36, y=9
        pixel_data[9][37] = 4'b0001; // x=37, y=9
        pixel_data[9][38] = 4'b0001; // x=38, y=9
        pixel_data[9][39] = 4'b0001; // x=39, y=9
        pixel_data[9][40] = 4'b0001; // x=40, y=9
        pixel_data[9][41] = 4'b0001; // x=41, y=9
        pixel_data[9][42] = 4'b0001; // x=42, y=9
        pixel_data[9][43] = 4'b0001; // x=43, y=9
        pixel_data[9][44] = 4'b0001; // x=44, y=9
        pixel_data[9][45] = 4'b0001; // x=45, y=9
        pixel_data[9][46] = 4'b0001; // x=46, y=9
        pixel_data[9][47] = 4'b0001; // x=47, y=9
        pixel_data[9][48] = 4'b0001; // x=48, y=9
        pixel_data[9][49] = 4'b0001; // x=49, y=9
        pixel_data[9][50] = 4'b0001; // x=50, y=9
        pixel_data[9][51] = 4'b0001; // x=51, y=9
        pixel_data[9][52] = 4'b0001; // x=52, y=9
        pixel_data[9][53] = 4'b0001; // x=53, y=9
        pixel_data[9][54] = 4'b0001; // x=54, y=9
        pixel_data[9][55] = 4'b0001; // x=55, y=9
        pixel_data[9][56] = 4'b0001; // x=56, y=9
        pixel_data[9][57] = 4'b0001; // x=57, y=9
        pixel_data[9][58] = 4'b0001; // x=58, y=9
        pixel_data[9][59] = 4'b0001; // x=59, y=9
        pixel_data[10][0] = 4'b0001; // x=0, y=10
        pixel_data[10][1] = 4'b0001; // x=1, y=10
        pixel_data[10][2] = 4'b0001; // x=2, y=10
        pixel_data[10][3] = 4'b0001; // x=3, y=10
        pixel_data[10][4] = 4'b0001; // x=4, y=10
        pixel_data[10][5] = 4'b0001; // x=5, y=10
        pixel_data[10][6] = 4'b0001; // x=6, y=10
        pixel_data[10][7] = 4'b0001; // x=7, y=10
        pixel_data[10][8] = 4'b0001; // x=8, y=10
        pixel_data[10][9] = 4'b0001; // x=9, y=10
        pixel_data[10][10] = 4'b0001; // x=10, y=10
        pixel_data[10][11] = 4'b0001; // x=11, y=10
        pixel_data[10][12] = 4'b0001; // x=12, y=10
        pixel_data[10][13] = 4'b0001; // x=13, y=10
        pixel_data[10][14] = 4'b0001; // x=14, y=10
        pixel_data[10][15] = 4'b0001; // x=15, y=10
        pixel_data[10][16] = 4'b0001; // x=16, y=10
        pixel_data[10][17] = 4'b0001; // x=17, y=10
        pixel_data[10][18] = 4'b0001; // x=18, y=10
        pixel_data[10][19] = 4'b0001; // x=19, y=10
        pixel_data[10][20] = 4'b0001; // x=20, y=10
        pixel_data[10][21] = 4'b0001; // x=21, y=10
        pixel_data[10][22] = 4'b0001; // x=22, y=10
        pixel_data[10][23] = 4'b0001; // x=23, y=10
        pixel_data[10][24] = 4'b0001; // x=24, y=10
        pixel_data[10][25] = 4'b0001; // x=25, y=10
        pixel_data[10][26] = 4'b0001; // x=26, y=10
        pixel_data[10][27] = 4'b0001; // x=27, y=10
        pixel_data[10][28] = 4'b0001; // x=28, y=10
        pixel_data[10][29] = 4'b0001; // x=29, y=10
        pixel_data[10][30] = 4'b0001; // x=30, y=10
        pixel_data[10][31] = 4'b0001; // x=31, y=10
        pixel_data[10][32] = 4'b0001; // x=32, y=10
        pixel_data[10][33] = 4'b0001; // x=33, y=10
        pixel_data[10][34] = 4'b0001; // x=34, y=10
        pixel_data[10][35] = 4'b0001; // x=35, y=10
        pixel_data[10][36] = 4'b0001; // x=36, y=10
        pixel_data[10][37] = 4'b0001; // x=37, y=10
        pixel_data[10][38] = 4'b0001; // x=38, y=10
        pixel_data[10][39] = 4'b0001; // x=39, y=10
        pixel_data[10][40] = 4'b0001; // x=40, y=10
        pixel_data[10][41] = 4'b0001; // x=41, y=10
        pixel_data[10][42] = 4'b0001; // x=42, y=10
        pixel_data[10][43] = 4'b0001; // x=43, y=10
        pixel_data[10][44] = 4'b0001; // x=44, y=10
        pixel_data[10][45] = 4'b0001; // x=45, y=10
        pixel_data[10][46] = 4'b0001; // x=46, y=10
        pixel_data[10][47] = 4'b0001; // x=47, y=10
        pixel_data[10][48] = 4'b0001; // x=48, y=10
        pixel_data[10][49] = 4'b0001; // x=49, y=10
        pixel_data[10][50] = 4'b0001; // x=50, y=10
        pixel_data[10][51] = 4'b0001; // x=51, y=10
        pixel_data[10][52] = 4'b0001; // x=52, y=10
        pixel_data[10][53] = 4'b0001; // x=53, y=10
        pixel_data[10][54] = 4'b0001; // x=54, y=10
        pixel_data[10][55] = 4'b0001; // x=55, y=10
        pixel_data[10][56] = 4'b0001; // x=56, y=10
        pixel_data[10][57] = 4'b0001; // x=57, y=10
        pixel_data[10][58] = 4'b0001; // x=58, y=10
        pixel_data[10][59] = 4'b0001; // x=59, y=10
        pixel_data[11][0] = 4'b0001; // x=0, y=11
        pixel_data[11][1] = 4'b0001; // x=1, y=11
        pixel_data[11][2] = 4'b0001; // x=2, y=11
        pixel_data[11][3] = 4'b0001; // x=3, y=11
        pixel_data[11][4] = 4'b0001; // x=4, y=11
        pixel_data[11][5] = 4'b0001; // x=5, y=11
        pixel_data[11][6] = 4'b0001; // x=6, y=11
        pixel_data[11][7] = 4'b0001; // x=7, y=11
        pixel_data[11][8] = 4'b0001; // x=8, y=11
        pixel_data[11][9] = 4'b0001; // x=9, y=11
        pixel_data[11][10] = 4'b0001; // x=10, y=11
        pixel_data[11][11] = 4'b0001; // x=11, y=11
        pixel_data[11][12] = 4'b0001; // x=12, y=11
        pixel_data[11][13] = 4'b0001; // x=13, y=11
        pixel_data[11][14] = 4'b0001; // x=14, y=11
        pixel_data[11][15] = 4'b0001; // x=15, y=11
        pixel_data[11][16] = 4'b0001; // x=16, y=11
        pixel_data[11][17] = 4'b0001; // x=17, y=11
        pixel_data[11][18] = 4'b0001; // x=18, y=11
        pixel_data[11][19] = 4'b0001; // x=19, y=11
        pixel_data[11][20] = 4'b0001; // x=20, y=11
        pixel_data[11][21] = 4'b0001; // x=21, y=11
        pixel_data[11][22] = 4'b0001; // x=22, y=11
        pixel_data[11][23] = 4'b0001; // x=23, y=11
        pixel_data[11][24] = 4'b0001; // x=24, y=11
        pixel_data[11][25] = 4'b0001; // x=25, y=11
        pixel_data[11][26] = 4'b0001; // x=26, y=11
        pixel_data[11][27] = 4'b0001; // x=27, y=11
        pixel_data[11][28] = 4'b0001; // x=28, y=11
        pixel_data[11][29] = 4'b0001; // x=29, y=11
        pixel_data[11][30] = 4'b0001; // x=30, y=11
        pixel_data[11][31] = 4'b0001; // x=31, y=11
        pixel_data[11][32] = 4'b0001; // x=32, y=11
        pixel_data[11][33] = 4'b0001; // x=33, y=11
        pixel_data[11][34] = 4'b0001; // x=34, y=11
        pixel_data[11][35] = 4'b0001; // x=35, y=11
        pixel_data[11][36] = 4'b0001; // x=36, y=11
        pixel_data[11][37] = 4'b0001; // x=37, y=11
        pixel_data[11][38] = 4'b0001; // x=38, y=11
        pixel_data[11][39] = 4'b0001; // x=39, y=11
        pixel_data[11][40] = 4'b0001; // x=40, y=11
        pixel_data[11][41] = 4'b0001; // x=41, y=11
        pixel_data[11][42] = 4'b0001; // x=42, y=11
        pixel_data[11][43] = 4'b0001; // x=43, y=11
        pixel_data[11][44] = 4'b0001; // x=44, y=11
        pixel_data[11][45] = 4'b0001; // x=45, y=11
        pixel_data[11][46] = 4'b0001; // x=46, y=11
        pixel_data[11][47] = 4'b0001; // x=47, y=11
        pixel_data[11][48] = 4'b0001; // x=48, y=11
        pixel_data[11][49] = 4'b0001; // x=49, y=11
        pixel_data[11][50] = 4'b0001; // x=50, y=11
        pixel_data[11][51] = 4'b0001; // x=51, y=11
        pixel_data[11][52] = 4'b0001; // x=52, y=11
        pixel_data[11][53] = 4'b0001; // x=53, y=11
        pixel_data[11][54] = 4'b0001; // x=54, y=11
        pixel_data[11][55] = 4'b0001; // x=55, y=11
        pixel_data[11][56] = 4'b0001; // x=56, y=11
        pixel_data[11][57] = 4'b0001; // x=57, y=11
        pixel_data[11][58] = 4'b0001; // x=58, y=11
        pixel_data[11][59] = 4'b0001; // x=59, y=11
        pixel_data[12][0] = 4'b0001; // x=0, y=12
        pixel_data[12][1] = 4'b0001; // x=1, y=12
        pixel_data[12][2] = 4'b0001; // x=2, y=12
        pixel_data[12][3] = 4'b0001; // x=3, y=12
        pixel_data[12][4] = 4'b0001; // x=4, y=12
        pixel_data[12][5] = 4'b0001; // x=5, y=12
        pixel_data[12][6] = 4'b0001; // x=6, y=12
        pixel_data[12][7] = 4'b0001; // x=7, y=12
        pixel_data[12][8] = 4'b0001; // x=8, y=12
        pixel_data[12][9] = 4'b0001; // x=9, y=12
        pixel_data[12][10] = 4'b0001; // x=10, y=12
        pixel_data[12][11] = 4'b0001; // x=11, y=12
        pixel_data[12][12] = 4'b0001; // x=12, y=12
        pixel_data[12][13] = 4'b0001; // x=13, y=12
        pixel_data[12][14] = 4'b0001; // x=14, y=12
        pixel_data[12][15] = 4'b0001; // x=15, y=12
        pixel_data[12][16] = 4'b0001; // x=16, y=12
        pixel_data[12][17] = 4'b0001; // x=17, y=12
        pixel_data[12][18] = 4'b0001; // x=18, y=12
        pixel_data[12][19] = 4'b0001; // x=19, y=12
        pixel_data[12][20] = 4'b0001; // x=20, y=12
        pixel_data[12][21] = 4'b0001; // x=21, y=12
        pixel_data[12][22] = 4'b0001; // x=22, y=12
        pixel_data[12][23] = 4'b0001; // x=23, y=12
        pixel_data[12][24] = 4'b0001; // x=24, y=12
        pixel_data[12][25] = 4'b0001; // x=25, y=12
        pixel_data[12][26] = 4'b0001; // x=26, y=12
        pixel_data[12][27] = 4'b0001; // x=27, y=12
        pixel_data[12][28] = 4'b0001; // x=28, y=12
        pixel_data[12][29] = 4'b0001; // x=29, y=12
        pixel_data[12][30] = 4'b0001; // x=30, y=12
        pixel_data[12][31] = 4'b0001; // x=31, y=12
        pixel_data[12][32] = 4'b0001; // x=32, y=12
        pixel_data[12][33] = 4'b0001; // x=33, y=12
        pixel_data[12][34] = 4'b0001; // x=34, y=12
        pixel_data[12][35] = 4'b0001; // x=35, y=12
        pixel_data[12][36] = 4'b0001; // x=36, y=12
        pixel_data[12][37] = 4'b0001; // x=37, y=12
        pixel_data[12][38] = 4'b0001; // x=38, y=12
        pixel_data[12][39] = 4'b0001; // x=39, y=12
        pixel_data[12][40] = 4'b0001; // x=40, y=12
        pixel_data[12][41] = 4'b0001; // x=41, y=12
        pixel_data[12][42] = 4'b0001; // x=42, y=12
        pixel_data[12][43] = 4'b0001; // x=43, y=12
        pixel_data[12][44] = 4'b0001; // x=44, y=12
        pixel_data[12][45] = 4'b0001; // x=45, y=12
        pixel_data[12][46] = 4'b0001; // x=46, y=12
        pixel_data[12][47] = 4'b0001; // x=47, y=12
        pixel_data[12][48] = 4'b0001; // x=48, y=12
        pixel_data[12][49] = 4'b0001; // x=49, y=12
        pixel_data[12][50] = 4'b0001; // x=50, y=12
        pixel_data[12][51] = 4'b0001; // x=51, y=12
        pixel_data[12][52] = 4'b0001; // x=52, y=12
        pixel_data[12][53] = 4'b0001; // x=53, y=12
        pixel_data[12][54] = 4'b0001; // x=54, y=12
        pixel_data[12][55] = 4'b0001; // x=55, y=12
        pixel_data[12][56] = 4'b0001; // x=56, y=12
        pixel_data[12][57] = 4'b0001; // x=57, y=12
        pixel_data[12][58] = 4'b0001; // x=58, y=12
        pixel_data[12][59] = 4'b0001; // x=59, y=12
        pixel_data[13][0] = 4'b0001; // x=0, y=13
        pixel_data[13][1] = 4'b0001; // x=1, y=13
        pixel_data[13][2] = 4'b0001; // x=2, y=13
        pixel_data[13][3] = 4'b0001; // x=3, y=13
        pixel_data[13][4] = 4'b0001; // x=4, y=13
        pixel_data[13][5] = 4'b0001; // x=5, y=13
        pixel_data[13][6] = 4'b0001; // x=6, y=13
        pixel_data[13][7] = 4'b0001; // x=7, y=13
        pixel_data[13][8] = 4'b0001; // x=8, y=13
        pixel_data[13][9] = 4'b0001; // x=9, y=13
        pixel_data[13][10] = 4'b0001; // x=10, y=13
        pixel_data[13][11] = 4'b0001; // x=11, y=13
        pixel_data[13][12] = 4'b0001; // x=12, y=13
        pixel_data[13][13] = 4'b0001; // x=13, y=13
        pixel_data[13][14] = 4'b0001; // x=14, y=13
        pixel_data[13][15] = 4'b0001; // x=15, y=13
        pixel_data[13][16] = 4'b0001; // x=16, y=13
        pixel_data[13][17] = 4'b0001; // x=17, y=13
        pixel_data[13][18] = 4'b0001; // x=18, y=13
        pixel_data[13][19] = 4'b0001; // x=19, y=13
        pixel_data[13][20] = 4'b0001; // x=20, y=13
        pixel_data[13][21] = 4'b0001; // x=21, y=13
        pixel_data[13][22] = 4'b0001; // x=22, y=13
        pixel_data[13][23] = 4'b0001; // x=23, y=13
        pixel_data[13][24] = 4'b0001; // x=24, y=13
        pixel_data[13][25] = 4'b0001; // x=25, y=13
        pixel_data[13][26] = 4'b0001; // x=26, y=13
        pixel_data[13][27] = 4'b0001; // x=27, y=13
        pixel_data[13][28] = 4'b0001; // x=28, y=13
        pixel_data[13][29] = 4'b0001; // x=29, y=13
        pixel_data[13][30] = 4'b0001; // x=30, y=13
        pixel_data[13][31] = 4'b0001; // x=31, y=13
        pixel_data[13][32] = 4'b0001; // x=32, y=13
        pixel_data[13][33] = 4'b0001; // x=33, y=13
        pixel_data[13][34] = 4'b0001; // x=34, y=13
        pixel_data[13][35] = 4'b0001; // x=35, y=13
        pixel_data[13][36] = 4'b0001; // x=36, y=13
        pixel_data[13][37] = 4'b0001; // x=37, y=13
        pixel_data[13][38] = 4'b0001; // x=38, y=13
        pixel_data[13][39] = 4'b0001; // x=39, y=13
        pixel_data[13][40] = 4'b0001; // x=40, y=13
        pixel_data[13][41] = 4'b0001; // x=41, y=13
        pixel_data[13][42] = 4'b0001; // x=42, y=13
        pixel_data[13][43] = 4'b0001; // x=43, y=13
        pixel_data[13][44] = 4'b0001; // x=44, y=13
        pixel_data[13][45] = 4'b0001; // x=45, y=13
        pixel_data[13][46] = 4'b0001; // x=46, y=13
        pixel_data[13][47] = 4'b0001; // x=47, y=13
        pixel_data[13][48] = 4'b0001; // x=48, y=13
        pixel_data[13][49] = 4'b0001; // x=49, y=13
        pixel_data[13][50] = 4'b0001; // x=50, y=13
        pixel_data[13][51] = 4'b0001; // x=51, y=13
        pixel_data[13][52] = 4'b0001; // x=52, y=13
        pixel_data[13][53] = 4'b0001; // x=53, y=13
        pixel_data[13][54] = 4'b0001; // x=54, y=13
        pixel_data[13][55] = 4'b0001; // x=55, y=13
        pixel_data[13][56] = 4'b0001; // x=56, y=13
        pixel_data[13][57] = 4'b0001; // x=57, y=13
        pixel_data[13][58] = 4'b0001; // x=58, y=13
        pixel_data[13][59] = 4'b0001; // x=59, y=13
        pixel_data[14][0] = 4'b0001; // x=0, y=14
        pixel_data[14][1] = 4'b0001; // x=1, y=14
        pixel_data[14][2] = 4'b0001; // x=2, y=14
        pixel_data[14][3] = 4'b0001; // x=3, y=14
        pixel_data[14][4] = 4'b0001; // x=4, y=14
        pixel_data[14][5] = 4'b0001; // x=5, y=14
        pixel_data[14][6] = 4'b0001; // x=6, y=14
        pixel_data[14][7] = 4'b0001; // x=7, y=14
        pixel_data[14][8] = 4'b0001; // x=8, y=14
        pixel_data[14][9] = 4'b0001; // x=9, y=14
        pixel_data[14][10] = 4'b0001; // x=10, y=14
        pixel_data[14][11] = 4'b0001; // x=11, y=14
        pixel_data[14][12] = 4'b0001; // x=12, y=14
        pixel_data[14][13] = 4'b0001; // x=13, y=14
        pixel_data[14][14] = 4'b0001; // x=14, y=14
        pixel_data[14][15] = 4'b0001; // x=15, y=14
        pixel_data[14][16] = 4'b0001; // x=16, y=14
        pixel_data[14][17] = 4'b0001; // x=17, y=14
        pixel_data[14][18] = 4'b0001; // x=18, y=14
        pixel_data[14][19] = 4'b0001; // x=19, y=14
        pixel_data[14][20] = 4'b0001; // x=20, y=14
        pixel_data[14][21] = 4'b0001; // x=21, y=14
        pixel_data[14][22] = 4'b0001; // x=22, y=14
        pixel_data[14][23] = 4'b0001; // x=23, y=14
        pixel_data[14][24] = 4'b0001; // x=24, y=14
        pixel_data[14][25] = 4'b0001; // x=25, y=14
        pixel_data[14][26] = 4'b0001; // x=26, y=14
        pixel_data[14][27] = 4'b0001; // x=27, y=14
        pixel_data[14][28] = 4'b0001; // x=28, y=14
        pixel_data[14][29] = 4'b0001; // x=29, y=14
        pixel_data[14][30] = 4'b0001; // x=30, y=14
        pixel_data[14][31] = 4'b0001; // x=31, y=14
        pixel_data[14][32] = 4'b0001; // x=32, y=14
        pixel_data[14][33] = 4'b0001; // x=33, y=14
        pixel_data[14][34] = 4'b0001; // x=34, y=14
        pixel_data[14][35] = 4'b0001; // x=35, y=14
        pixel_data[14][36] = 4'b0001; // x=36, y=14
        pixel_data[14][37] = 4'b0001; // x=37, y=14
        pixel_data[14][38] = 4'b0001; // x=38, y=14
        pixel_data[14][39] = 4'b0001; // x=39, y=14
        pixel_data[14][40] = 4'b0001; // x=40, y=14
        pixel_data[14][41] = 4'b0001; // x=41, y=14
        pixel_data[14][42] = 4'b0001; // x=42, y=14
        pixel_data[14][43] = 4'b0001; // x=43, y=14
        pixel_data[14][44] = 4'b0001; // x=44, y=14
        pixel_data[14][45] = 4'b0001; // x=45, y=14
        pixel_data[14][46] = 4'b0001; // x=46, y=14
        pixel_data[14][47] = 4'b0001; // x=47, y=14
        pixel_data[14][48] = 4'b0001; // x=48, y=14
        pixel_data[14][49] = 4'b0001; // x=49, y=14
        pixel_data[14][50] = 4'b0001; // x=50, y=14
        pixel_data[14][51] = 4'b0001; // x=51, y=14
        pixel_data[14][52] = 4'b0001; // x=52, y=14
        pixel_data[14][53] = 4'b0001; // x=53, y=14
        pixel_data[14][54] = 4'b0001; // x=54, y=14
        pixel_data[14][55] = 4'b0001; // x=55, y=14
        pixel_data[14][56] = 4'b0001; // x=56, y=14
        pixel_data[14][57] = 4'b0001; // x=57, y=14
        pixel_data[14][58] = 4'b0001; // x=58, y=14
        pixel_data[14][59] = 4'b0001; // x=59, y=14
        pixel_data[15][0] = 4'b0001; // x=0, y=15
        pixel_data[15][1] = 4'b0001; // x=1, y=15
        pixel_data[15][2] = 4'b0001; // x=2, y=15
        pixel_data[15][3] = 4'b0001; // x=3, y=15
        pixel_data[15][4] = 4'b0001; // x=4, y=15
        pixel_data[15][5] = 4'b0001; // x=5, y=15
        pixel_data[15][6] = 4'b0001; // x=6, y=15
        pixel_data[15][7] = 4'b0001; // x=7, y=15
        pixel_data[15][8] = 4'b0001; // x=8, y=15
        pixel_data[15][9] = 4'b0001; // x=9, y=15
        pixel_data[15][10] = 4'b0001; // x=10, y=15
        pixel_data[15][11] = 4'b0001; // x=11, y=15
        pixel_data[15][12] = 4'b0001; // x=12, y=15
        pixel_data[15][13] = 4'b0001; // x=13, y=15
        pixel_data[15][14] = 4'b0001; // x=14, y=15
        pixel_data[15][15] = 4'b0001; // x=15, y=15
        pixel_data[15][16] = 4'b0001; // x=16, y=15
        pixel_data[15][17] = 4'b0001; // x=17, y=15
        pixel_data[15][18] = 4'b0001; // x=18, y=15
        pixel_data[15][19] = 4'b0001; // x=19, y=15
        pixel_data[15][20] = 4'b0001; // x=20, y=15
        pixel_data[15][21] = 4'b0001; // x=21, y=15
        pixel_data[15][22] = 4'b0001; // x=22, y=15
        pixel_data[15][23] = 4'b0001; // x=23, y=15
        pixel_data[15][24] = 4'b0001; // x=24, y=15
        pixel_data[15][25] = 4'b0001; // x=25, y=15
        pixel_data[15][26] = 4'b0001; // x=26, y=15
        pixel_data[15][27] = 4'b0001; // x=27, y=15
        pixel_data[15][28] = 4'b0001; // x=28, y=15
        pixel_data[15][29] = 4'b0001; // x=29, y=15
        pixel_data[15][30] = 4'b0001; // x=30, y=15
        pixel_data[15][31] = 4'b0001; // x=31, y=15
        pixel_data[15][32] = 4'b0001; // x=32, y=15
        pixel_data[15][33] = 4'b0001; // x=33, y=15
        pixel_data[15][34] = 4'b0001; // x=34, y=15
        pixel_data[15][35] = 4'b0001; // x=35, y=15
        pixel_data[15][36] = 4'b0001; // x=36, y=15
        pixel_data[15][37] = 4'b0001; // x=37, y=15
        pixel_data[15][38] = 4'b0001; // x=38, y=15
        pixel_data[15][39] = 4'b0001; // x=39, y=15
        pixel_data[15][40] = 4'b0001; // x=40, y=15
        pixel_data[15][41] = 4'b0001; // x=41, y=15
        pixel_data[15][42] = 4'b0001; // x=42, y=15
        pixel_data[15][43] = 4'b0001; // x=43, y=15
        pixel_data[15][44] = 4'b0001; // x=44, y=15
        pixel_data[15][45] = 4'b0001; // x=45, y=15
        pixel_data[15][46] = 4'b0001; // x=46, y=15
        pixel_data[15][47] = 4'b0001; // x=47, y=15
        pixel_data[15][48] = 4'b0001; // x=48, y=15
        pixel_data[15][49] = 4'b0001; // x=49, y=15
        pixel_data[15][50] = 4'b0001; // x=50, y=15
        pixel_data[15][51] = 4'b0001; // x=51, y=15
        pixel_data[15][52] = 4'b0001; // x=52, y=15
        pixel_data[15][53] = 4'b0001; // x=53, y=15
        pixel_data[15][54] = 4'b0001; // x=54, y=15
        pixel_data[15][55] = 4'b0001; // x=55, y=15
        pixel_data[15][56] = 4'b0001; // x=56, y=15
        pixel_data[15][57] = 4'b0001; // x=57, y=15
        pixel_data[15][58] = 4'b0001; // x=58, y=15
        pixel_data[15][59] = 4'b0001; // x=59, y=15
        pixel_data[16][0] = 4'b0001; // x=0, y=16
        pixel_data[16][1] = 4'b0001; // x=1, y=16
        pixel_data[16][2] = 4'b0001; // x=2, y=16
        pixel_data[16][3] = 4'b0001; // x=3, y=16
        pixel_data[16][4] = 4'b0001; // x=4, y=16
        pixel_data[16][5] = 4'b0001; // x=5, y=16
        pixel_data[16][6] = 4'b0001; // x=6, y=16
        pixel_data[16][7] = 4'b0001; // x=7, y=16
        pixel_data[16][8] = 4'b0001; // x=8, y=16
        pixel_data[16][9] = 4'b0001; // x=9, y=16
        pixel_data[16][10] = 4'b0001; // x=10, y=16
        pixel_data[16][11] = 4'b0001; // x=11, y=16
        pixel_data[16][12] = 4'b0001; // x=12, y=16
        pixel_data[16][13] = 4'b0001; // x=13, y=16
        pixel_data[16][14] = 4'b0001; // x=14, y=16
        pixel_data[16][15] = 4'b0001; // x=15, y=16
        pixel_data[16][16] = 4'b0001; // x=16, y=16
        pixel_data[16][17] = 4'b0001; // x=17, y=16
        pixel_data[16][18] = 4'b0001; // x=18, y=16
        pixel_data[16][19] = 4'b0001; // x=19, y=16
        pixel_data[16][20] = 4'b0001; // x=20, y=16
        pixel_data[16][21] = 4'b0001; // x=21, y=16
        pixel_data[16][22] = 4'b0001; // x=22, y=16
        pixel_data[16][23] = 4'b0001; // x=23, y=16
        pixel_data[16][24] = 4'b0001; // x=24, y=16
        pixel_data[16][25] = 4'b0001; // x=25, y=16
        pixel_data[16][26] = 4'b0001; // x=26, y=16
        pixel_data[16][27] = 4'b0001; // x=27, y=16
        pixel_data[16][28] = 4'b0001; // x=28, y=16
        pixel_data[16][29] = 4'b0001; // x=29, y=16
        pixel_data[16][30] = 4'b0001; // x=30, y=16
        pixel_data[16][31] = 4'b0001; // x=31, y=16
        pixel_data[16][32] = 4'b0001; // x=32, y=16
        pixel_data[16][33] = 4'b0001; // x=33, y=16
        pixel_data[16][34] = 4'b0001; // x=34, y=16
        pixel_data[16][35] = 4'b0001; // x=35, y=16
        pixel_data[16][36] = 4'b0001; // x=36, y=16
        pixel_data[16][37] = 4'b0001; // x=37, y=16
        pixel_data[16][38] = 4'b0001; // x=38, y=16
        pixel_data[16][39] = 4'b0001; // x=39, y=16
        pixel_data[16][40] = 4'b0001; // x=40, y=16
        pixel_data[16][41] = 4'b0001; // x=41, y=16
        pixel_data[16][42] = 4'b0001; // x=42, y=16
        pixel_data[16][43] = 4'b0001; // x=43, y=16
        pixel_data[16][44] = 4'b0001; // x=44, y=16
        pixel_data[16][45] = 4'b0001; // x=45, y=16
        pixel_data[16][46] = 4'b0001; // x=46, y=16
        pixel_data[16][47] = 4'b0001; // x=47, y=16
        pixel_data[16][48] = 4'b0001; // x=48, y=16
        pixel_data[16][49] = 4'b0001; // x=49, y=16
        pixel_data[16][50] = 4'b0001; // x=50, y=16
        pixel_data[16][51] = 4'b0001; // x=51, y=16
        pixel_data[16][52] = 4'b0001; // x=52, y=16
        pixel_data[16][53] = 4'b0001; // x=53, y=16
        pixel_data[16][54] = 4'b0001; // x=54, y=16
        pixel_data[16][55] = 4'b0001; // x=55, y=16
        pixel_data[16][56] = 4'b0001; // x=56, y=16
        pixel_data[16][57] = 4'b0001; // x=57, y=16
        pixel_data[16][58] = 4'b0001; // x=58, y=16
        pixel_data[16][59] = 4'b0001; // x=59, y=16
        pixel_data[17][0] = 4'b0001; // x=0, y=17
        pixel_data[17][1] = 4'b0001; // x=1, y=17
        pixel_data[17][2] = 4'b0001; // x=2, y=17
        pixel_data[17][3] = 4'b0001; // x=3, y=17
        pixel_data[17][4] = 4'b0001; // x=4, y=17
        pixel_data[17][5] = 4'b0001; // x=5, y=17
        pixel_data[17][6] = 4'b0001; // x=6, y=17
        pixel_data[17][7] = 4'b0001; // x=7, y=17
        pixel_data[17][8] = 4'b0001; // x=8, y=17
        pixel_data[17][9] = 4'b0001; // x=9, y=17
        pixel_data[17][10] = 4'b0001; // x=10, y=17
        pixel_data[17][11] = 4'b0001; // x=11, y=17
        pixel_data[17][12] = 4'b0001; // x=12, y=17
        pixel_data[17][13] = 4'b0001; // x=13, y=17
        pixel_data[17][14] = 4'b0001; // x=14, y=17
        pixel_data[17][15] = 4'b1011; // x=15, y=17
        pixel_data[17][16] = 4'b1011; // x=16, y=17
        pixel_data[17][17] = 4'b1000; // x=17, y=17
        pixel_data[17][18] = 4'b1000; // x=18, y=17
        pixel_data[17][19] = 4'b1000; // x=19, y=17
        pixel_data[17][20] = 4'b1000; // x=20, y=17
        pixel_data[17][21] = 4'b1000; // x=21, y=17
        pixel_data[17][22] = 4'b1000; // x=22, y=17
        pixel_data[17][23] = 4'b1000; // x=23, y=17
        pixel_data[17][24] = 4'b1000; // x=24, y=17
        pixel_data[17][25] = 4'b1000; // x=25, y=17
        pixel_data[17][26] = 4'b1000; // x=26, y=17
        pixel_data[17][27] = 4'b1000; // x=27, y=17
        pixel_data[17][28] = 4'b1000; // x=28, y=17
        pixel_data[17][29] = 4'b1000; // x=29, y=17
        pixel_data[17][30] = 4'b1000; // x=30, y=17
        pixel_data[17][31] = 4'b1000; // x=31, y=17
        pixel_data[17][32] = 4'b1000; // x=32, y=17
        pixel_data[17][33] = 4'b1000; // x=33, y=17
        pixel_data[17][34] = 4'b1000; // x=34, y=17
        pixel_data[17][35] = 4'b1000; // x=35, y=17
        pixel_data[17][36] = 4'b1000; // x=36, y=17
        pixel_data[17][37] = 4'b1000; // x=37, y=17
        pixel_data[17][38] = 4'b1000; // x=38, y=17
        pixel_data[17][39] = 4'b1000; // x=39, y=17
        pixel_data[17][40] = 4'b1011; // x=40, y=17
        pixel_data[17][41] = 4'b0001; // x=41, y=17
        pixel_data[17][42] = 4'b0001; // x=42, y=17
        pixel_data[17][43] = 4'b0001; // x=43, y=17
        pixel_data[17][44] = 4'b0001; // x=44, y=17
        pixel_data[17][45] = 4'b0001; // x=45, y=17
        pixel_data[17][46] = 4'b0001; // x=46, y=17
        pixel_data[17][47] = 4'b0001; // x=47, y=17
        pixel_data[17][48] = 4'b0001; // x=48, y=17
        pixel_data[17][49] = 4'b0001; // x=49, y=17
        pixel_data[17][50] = 4'b0001; // x=50, y=17
        pixel_data[17][51] = 4'b0001; // x=51, y=17
        pixel_data[17][52] = 4'b0001; // x=52, y=17
        pixel_data[17][53] = 4'b0001; // x=53, y=17
        pixel_data[17][54] = 4'b0001; // x=54, y=17
        pixel_data[17][55] = 4'b0001; // x=55, y=17
        pixel_data[17][56] = 4'b0001; // x=56, y=17
        pixel_data[17][57] = 4'b0001; // x=57, y=17
        pixel_data[17][58] = 4'b0001; // x=58, y=17
        pixel_data[17][59] = 4'b0001; // x=59, y=17
        pixel_data[18][0] = 4'b0001; // x=0, y=18
        pixel_data[18][1] = 4'b0001; // x=1, y=18
        pixel_data[18][2] = 4'b0001; // x=2, y=18
        pixel_data[18][3] = 4'b0001; // x=3, y=18
        pixel_data[18][4] = 4'b0001; // x=4, y=18
        pixel_data[18][5] = 4'b0001; // x=5, y=18
        pixel_data[18][6] = 4'b0001; // x=6, y=18
        pixel_data[18][7] = 4'b0001; // x=7, y=18
        pixel_data[18][8] = 4'b0001; // x=8, y=18
        pixel_data[18][9] = 4'b0001; // x=9, y=18
        pixel_data[18][10] = 4'b0001; // x=10, y=18
        pixel_data[18][11] = 4'b0001; // x=11, y=18
        pixel_data[18][12] = 4'b0001; // x=12, y=18
        pixel_data[18][13] = 4'b0001; // x=13, y=18
        pixel_data[18][14] = 4'b1011; // x=14, y=18
        pixel_data[18][15] = 4'b0001; // x=15, y=18
        pixel_data[18][16] = 4'b0011; // x=16, y=18
        pixel_data[18][17] = 4'b0100; // x=17, y=18
        pixel_data[18][18] = 4'b0100; // x=18, y=18
        pixel_data[18][19] = 4'b0100; // x=19, y=18
        pixel_data[18][20] = 4'b0100; // x=20, y=18
        pixel_data[18][21] = 4'b0100; // x=21, y=18
        pixel_data[18][22] = 4'b0100; // x=22, y=18
        pixel_data[18][23] = 4'b0100; // x=23, y=18
        pixel_data[18][24] = 4'b0100; // x=24, y=18
        pixel_data[18][25] = 4'b0100; // x=25, y=18
        pixel_data[18][26] = 4'b0100; // x=26, y=18
        pixel_data[18][27] = 4'b0100; // x=27, y=18
        pixel_data[18][28] = 4'b0100; // x=28, y=18
        pixel_data[18][29] = 4'b0100; // x=29, y=18
        pixel_data[18][30] = 4'b0100; // x=30, y=18
        pixel_data[18][31] = 4'b0100; // x=31, y=18
        pixel_data[18][32] = 4'b0100; // x=32, y=18
        pixel_data[18][33] = 4'b0100; // x=33, y=18
        pixel_data[18][34] = 4'b0100; // x=34, y=18
        pixel_data[18][35] = 4'b0100; // x=35, y=18
        pixel_data[18][36] = 4'b0100; // x=36, y=18
        pixel_data[18][37] = 4'b0100; // x=37, y=18
        pixel_data[18][38] = 4'b0100; // x=38, y=18
        pixel_data[18][39] = 4'b0100; // x=39, y=18
        pixel_data[18][40] = 4'b0111; // x=40, y=18
        pixel_data[18][41] = 4'b1000; // x=41, y=18
        pixel_data[18][42] = 4'b0001; // x=42, y=18
        pixel_data[18][43] = 4'b0001; // x=43, y=18
        pixel_data[18][44] = 4'b0001; // x=44, y=18
        pixel_data[18][45] = 4'b0001; // x=45, y=18
        pixel_data[18][46] = 4'b0001; // x=46, y=18
        pixel_data[18][47] = 4'b0001; // x=47, y=18
        pixel_data[18][48] = 4'b0001; // x=48, y=18
        pixel_data[18][49] = 4'b0001; // x=49, y=18
        pixel_data[18][50] = 4'b0001; // x=50, y=18
        pixel_data[18][51] = 4'b0001; // x=51, y=18
        pixel_data[18][52] = 4'b0001; // x=52, y=18
        pixel_data[18][53] = 4'b0001; // x=53, y=18
        pixel_data[18][54] = 4'b0001; // x=54, y=18
        pixel_data[18][55] = 4'b0001; // x=55, y=18
        pixel_data[18][56] = 4'b0001; // x=56, y=18
        pixel_data[18][57] = 4'b0001; // x=57, y=18
        pixel_data[18][58] = 4'b0001; // x=58, y=18
        pixel_data[18][59] = 4'b0001; // x=59, y=18
        pixel_data[19][0] = 4'b0001; // x=0, y=19
        pixel_data[19][1] = 4'b0001; // x=1, y=19
        pixel_data[19][2] = 4'b0001; // x=2, y=19
        pixel_data[19][3] = 4'b0001; // x=3, y=19
        pixel_data[19][4] = 4'b0001; // x=4, y=19
        pixel_data[19][5] = 4'b0001; // x=5, y=19
        pixel_data[19][6] = 4'b0001; // x=6, y=19
        pixel_data[19][7] = 4'b0001; // x=7, y=19
        pixel_data[19][8] = 4'b0001; // x=8, y=19
        pixel_data[19][9] = 4'b0001; // x=9, y=19
        pixel_data[19][10] = 4'b0001; // x=10, y=19
        pixel_data[19][11] = 4'b0001; // x=11, y=19
        pixel_data[19][12] = 4'b0001; // x=12, y=19
        pixel_data[19][13] = 4'b0001; // x=13, y=19
        pixel_data[19][14] = 4'b1011; // x=14, y=19
        pixel_data[19][15] = 4'b0001; // x=15, y=19
        pixel_data[19][16] = 4'b1001; // x=16, y=19
        pixel_data[19][17] = 4'b1010; // x=17, y=19
        pixel_data[19][18] = 4'b1010; // x=18, y=19
        pixel_data[19][19] = 4'b1010; // x=19, y=19
        pixel_data[19][20] = 4'b1010; // x=20, y=19
        pixel_data[19][21] = 4'b1010; // x=21, y=19
        pixel_data[19][22] = 4'b1010; // x=22, y=19
        pixel_data[19][23] = 4'b1010; // x=23, y=19
        pixel_data[19][24] = 4'b1010; // x=24, y=19
        pixel_data[19][25] = 4'b1010; // x=25, y=19
        pixel_data[19][26] = 4'b1010; // x=26, y=19
        pixel_data[19][27] = 4'b1010; // x=27, y=19
        pixel_data[19][28] = 4'b1010; // x=28, y=19
        pixel_data[19][29] = 4'b1010; // x=29, y=19
        pixel_data[19][30] = 4'b1010; // x=30, y=19
        pixel_data[19][31] = 4'b1010; // x=31, y=19
        pixel_data[19][32] = 4'b1010; // x=32, y=19
        pixel_data[19][33] = 4'b1010; // x=33, y=19
        pixel_data[19][34] = 4'b1010; // x=34, y=19
        pixel_data[19][35] = 4'b1010; // x=35, y=19
        pixel_data[19][36] = 4'b1010; // x=36, y=19
        pixel_data[19][37] = 4'b1010; // x=37, y=19
        pixel_data[19][38] = 4'b1010; // x=38, y=19
        pixel_data[19][39] = 4'b1010; // x=39, y=19
        pixel_data[19][40] = 4'b1010; // x=40, y=19
        pixel_data[19][41] = 4'b0110; // x=41, y=19
        pixel_data[19][42] = 4'b0001; // x=42, y=19
        pixel_data[19][43] = 4'b1011; // x=43, y=19
        pixel_data[19][44] = 4'b0001; // x=44, y=19
        pixel_data[19][45] = 4'b0001; // x=45, y=19
        pixel_data[19][46] = 4'b0001; // x=46, y=19
        pixel_data[19][47] = 4'b0001; // x=47, y=19
        pixel_data[19][48] = 4'b0001; // x=48, y=19
        pixel_data[19][49] = 4'b0001; // x=49, y=19
        pixel_data[19][50] = 4'b0001; // x=50, y=19
        pixel_data[19][51] = 4'b0001; // x=51, y=19
        pixel_data[19][52] = 4'b0001; // x=52, y=19
        pixel_data[19][53] = 4'b0001; // x=53, y=19
        pixel_data[19][54] = 4'b0001; // x=54, y=19
        pixel_data[19][55] = 4'b0001; // x=55, y=19
        pixel_data[19][56] = 4'b0001; // x=56, y=19
        pixel_data[19][57] = 4'b0001; // x=57, y=19
        pixel_data[19][58] = 4'b0001; // x=58, y=19
        pixel_data[19][59] = 4'b0001; // x=59, y=19
        pixel_data[20][0] = 4'b0001; // x=0, y=20
        pixel_data[20][1] = 4'b0001; // x=1, y=20
        pixel_data[20][2] = 4'b0001; // x=2, y=20
        pixel_data[20][3] = 4'b0001; // x=3, y=20
        pixel_data[20][4] = 4'b0001; // x=4, y=20
        pixel_data[20][5] = 4'b0001; // x=5, y=20
        pixel_data[20][6] = 4'b0001; // x=6, y=20
        pixel_data[20][7] = 4'b0001; // x=7, y=20
        pixel_data[20][8] = 4'b0001; // x=8, y=20
        pixel_data[20][9] = 4'b0001; // x=9, y=20
        pixel_data[20][10] = 4'b0001; // x=10, y=20
        pixel_data[20][11] = 4'b0001; // x=11, y=20
        pixel_data[20][12] = 4'b0001; // x=12, y=20
        pixel_data[20][13] = 4'b0001; // x=13, y=20
        pixel_data[20][14] = 4'b1011; // x=14, y=20
        pixel_data[20][15] = 4'b0001; // x=15, y=20
        pixel_data[20][16] = 4'b0011; // x=16, y=20
        pixel_data[20][17] = 4'b0010; // x=17, y=20
        pixel_data[20][18] = 4'b0010; // x=18, y=20
        pixel_data[20][19] = 4'b0010; // x=19, y=20
        pixel_data[20][20] = 4'b0010; // x=20, y=20
        pixel_data[20][21] = 4'b0010; // x=21, y=20
        pixel_data[20][22] = 4'b0010; // x=22, y=20
        pixel_data[20][23] = 4'b0010; // x=23, y=20
        pixel_data[20][24] = 4'b0010; // x=24, y=20
        pixel_data[20][25] = 4'b0010; // x=25, y=20
        pixel_data[20][26] = 4'b0010; // x=26, y=20
        pixel_data[20][27] = 4'b0010; // x=27, y=20
        pixel_data[20][28] = 4'b0010; // x=28, y=20
        pixel_data[20][29] = 4'b0010; // x=29, y=20
        pixel_data[20][30] = 4'b0010; // x=30, y=20
        pixel_data[20][31] = 4'b0010; // x=31, y=20
        pixel_data[20][32] = 4'b0010; // x=32, y=20
        pixel_data[20][33] = 4'b0010; // x=33, y=20
        pixel_data[20][34] = 4'b1010; // x=34, y=20
        pixel_data[20][35] = 4'b1010; // x=35, y=20
        pixel_data[20][36] = 4'b1010; // x=36, y=20
        pixel_data[20][37] = 4'b0010; // x=37, y=20
        pixel_data[20][38] = 4'b0010; // x=38, y=20
        pixel_data[20][39] = 4'b0010; // x=39, y=20
        pixel_data[20][40] = 4'b1010; // x=40, y=20
        pixel_data[20][41] = 4'b1100; // x=41, y=20
        pixel_data[20][42] = 4'b0001; // x=42, y=20
        pixel_data[20][43] = 4'b1011; // x=43, y=20
        pixel_data[20][44] = 4'b0001; // x=44, y=20
        pixel_data[20][45] = 4'b0001; // x=45, y=20
        pixel_data[20][46] = 4'b0001; // x=46, y=20
        pixel_data[20][47] = 4'b0001; // x=47, y=20
        pixel_data[20][48] = 4'b0001; // x=48, y=20
        pixel_data[20][49] = 4'b0001; // x=49, y=20
        pixel_data[20][50] = 4'b0001; // x=50, y=20
        pixel_data[20][51] = 4'b0001; // x=51, y=20
        pixel_data[20][52] = 4'b0001; // x=52, y=20
        pixel_data[20][53] = 4'b0001; // x=53, y=20
        pixel_data[20][54] = 4'b0001; // x=54, y=20
        pixel_data[20][55] = 4'b0001; // x=55, y=20
        pixel_data[20][56] = 4'b0001; // x=56, y=20
        pixel_data[20][57] = 4'b0001; // x=57, y=20
        pixel_data[20][58] = 4'b0001; // x=58, y=20
        pixel_data[20][59] = 4'b0001; // x=59, y=20
        pixel_data[21][0] = 4'b0001; // x=0, y=21
        pixel_data[21][1] = 4'b0001; // x=1, y=21
        pixel_data[21][2] = 4'b0001; // x=2, y=21
        pixel_data[21][3] = 4'b0001; // x=3, y=21
        pixel_data[21][4] = 4'b0001; // x=4, y=21
        pixel_data[21][5] = 4'b0001; // x=5, y=21
        pixel_data[21][6] = 4'b0001; // x=6, y=21
        pixel_data[21][7] = 4'b0001; // x=7, y=21
        pixel_data[21][8] = 4'b0001; // x=8, y=21
        pixel_data[21][9] = 4'b0001; // x=9, y=21
        pixel_data[21][10] = 4'b0001; // x=10, y=21
        pixel_data[21][11] = 4'b0001; // x=11, y=21
        pixel_data[21][12] = 4'b0001; // x=12, y=21
        pixel_data[21][13] = 4'b0001; // x=13, y=21
        pixel_data[21][14] = 4'b1011; // x=14, y=21
        pixel_data[21][15] = 4'b0001; // x=15, y=21
        pixel_data[21][16] = 4'b1001; // x=16, y=21
        pixel_data[21][17] = 4'b1010; // x=17, y=21
        pixel_data[21][18] = 4'b1010; // x=18, y=21
        pixel_data[21][19] = 4'b1010; // x=19, y=21
        pixel_data[21][20] = 4'b1010; // x=20, y=21
        pixel_data[21][21] = 4'b1010; // x=21, y=21
        pixel_data[21][22] = 4'b1010; // x=22, y=21
        pixel_data[21][23] = 4'b1010; // x=23, y=21
        pixel_data[21][24] = 4'b1010; // x=24, y=21
        pixel_data[21][25] = 4'b1010; // x=25, y=21
        pixel_data[21][26] = 4'b1010; // x=26, y=21
        pixel_data[21][27] = 4'b1010; // x=27, y=21
        pixel_data[21][28] = 4'b1010; // x=28, y=21
        pixel_data[21][29] = 4'b1010; // x=29, y=21
        pixel_data[21][30] = 4'b1010; // x=30, y=21
        pixel_data[21][31] = 4'b1010; // x=31, y=21
        pixel_data[21][32] = 4'b1010; // x=32, y=21
        pixel_data[21][33] = 4'b1010; // x=33, y=21
        pixel_data[21][34] = 4'b1010; // x=34, y=21
        pixel_data[21][35] = 4'b1010; // x=35, y=21
        pixel_data[21][36] = 4'b0010; // x=36, y=21
        pixel_data[21][37] = 4'b0010; // x=37, y=21
        pixel_data[21][38] = 4'b1010; // x=38, y=21
        pixel_data[21][39] = 4'b0010; // x=39, y=21
        pixel_data[21][40] = 4'b0010; // x=40, y=21
        pixel_data[21][41] = 4'b0011; // x=41, y=21
        pixel_data[21][42] = 4'b0001; // x=42, y=21
        pixel_data[21][43] = 4'b0001; // x=43, y=21
        pixel_data[21][44] = 4'b0001; // x=44, y=21
        pixel_data[21][45] = 4'b0001; // x=45, y=21
        pixel_data[21][46] = 4'b0001; // x=46, y=21
        pixel_data[21][47] = 4'b0001; // x=47, y=21
        pixel_data[21][48] = 4'b0001; // x=48, y=21
        pixel_data[21][49] = 4'b0001; // x=49, y=21
        pixel_data[21][50] = 4'b0001; // x=50, y=21
        pixel_data[21][51] = 4'b0001; // x=51, y=21
        pixel_data[21][52] = 4'b0001; // x=52, y=21
        pixel_data[21][53] = 4'b0001; // x=53, y=21
        pixel_data[21][54] = 4'b0001; // x=54, y=21
        pixel_data[21][55] = 4'b0001; // x=55, y=21
        pixel_data[21][56] = 4'b0001; // x=56, y=21
        pixel_data[21][57] = 4'b0001; // x=57, y=21
        pixel_data[21][58] = 4'b0001; // x=58, y=21
        pixel_data[21][59] = 4'b0001; // x=59, y=21
        pixel_data[22][0] = 4'b0001; // x=0, y=22
        pixel_data[22][1] = 4'b0001; // x=1, y=22
        pixel_data[22][2] = 4'b0001; // x=2, y=22
        pixel_data[22][3] = 4'b0001; // x=3, y=22
        pixel_data[22][4] = 4'b0001; // x=4, y=22
        pixel_data[22][5] = 4'b0001; // x=5, y=22
        pixel_data[22][6] = 4'b0001; // x=6, y=22
        pixel_data[22][7] = 4'b0001; // x=7, y=22
        pixel_data[22][8] = 4'b0001; // x=8, y=22
        pixel_data[22][9] = 4'b0001; // x=9, y=22
        pixel_data[22][10] = 4'b0001; // x=10, y=22
        pixel_data[22][11] = 4'b0001; // x=11, y=22
        pixel_data[22][12] = 4'b0001; // x=12, y=22
        pixel_data[22][13] = 4'b0001; // x=13, y=22
        pixel_data[22][14] = 4'b1011; // x=14, y=22
        pixel_data[22][15] = 4'b0001; // x=15, y=22
        pixel_data[22][16] = 4'b1111; // x=16, y=22
        pixel_data[22][17] = 4'b0000; // x=17, y=22
        pixel_data[22][18] = 4'b0000; // x=18, y=22
        pixel_data[22][19] = 4'b0000; // x=19, y=22
        pixel_data[22][20] = 4'b0000; // x=20, y=22
        pixel_data[22][21] = 4'b0000; // x=21, y=22
        pixel_data[22][22] = 4'b0000; // x=22, y=22
        pixel_data[22][23] = 4'b0000; // x=23, y=22
        pixel_data[22][24] = 4'b0000; // x=24, y=22
        pixel_data[22][25] = 4'b0000; // x=25, y=22
        pixel_data[22][26] = 4'b0000; // x=26, y=22
        pixel_data[22][27] = 4'b0000; // x=27, y=22
        pixel_data[22][28] = 4'b0000; // x=28, y=22
        pixel_data[22][29] = 4'b0000; // x=29, y=22
        pixel_data[22][30] = 4'b0000; // x=30, y=22
        pixel_data[22][31] = 4'b0000; // x=31, y=22
        pixel_data[22][32] = 4'b0000; // x=32, y=22
        pixel_data[22][33] = 4'b0100; // x=33, y=22
        pixel_data[22][34] = 4'b1010; // x=34, y=22
        pixel_data[22][35] = 4'b0010; // x=35, y=22
        pixel_data[22][36] = 4'b1010; // x=36, y=22
        pixel_data[22][37] = 4'b0010; // x=37, y=22
        pixel_data[22][38] = 4'b0010; // x=38, y=22
        pixel_data[22][39] = 4'b1010; // x=39, y=22
        pixel_data[22][40] = 4'b1101; // x=40, y=22
        pixel_data[22][41] = 4'b0001; // x=41, y=22
        pixel_data[22][42] = 4'b1011; // x=42, y=22
        pixel_data[22][43] = 4'b0001; // x=43, y=22
        pixel_data[22][44] = 4'b0001; // x=44, y=22
        pixel_data[22][45] = 4'b0001; // x=45, y=22
        pixel_data[22][46] = 4'b0001; // x=46, y=22
        pixel_data[22][47] = 4'b0001; // x=47, y=22
        pixel_data[22][48] = 4'b0001; // x=48, y=22
        pixel_data[22][49] = 4'b0001; // x=49, y=22
        pixel_data[22][50] = 4'b0001; // x=50, y=22
        pixel_data[22][51] = 4'b0001; // x=51, y=22
        pixel_data[22][52] = 4'b0001; // x=52, y=22
        pixel_data[22][53] = 4'b0001; // x=53, y=22
        pixel_data[22][54] = 4'b0001; // x=54, y=22
        pixel_data[22][55] = 4'b0001; // x=55, y=22
        pixel_data[22][56] = 4'b0001; // x=56, y=22
        pixel_data[22][57] = 4'b0001; // x=57, y=22
        pixel_data[22][58] = 4'b0001; // x=58, y=22
        pixel_data[22][59] = 4'b0001; // x=59, y=22
        pixel_data[23][0] = 4'b0001; // x=0, y=23
        pixel_data[23][1] = 4'b0001; // x=1, y=23
        pixel_data[23][2] = 4'b0001; // x=2, y=23
        pixel_data[23][3] = 4'b0001; // x=3, y=23
        pixel_data[23][4] = 4'b0001; // x=4, y=23
        pixel_data[23][5] = 4'b0001; // x=5, y=23
        pixel_data[23][6] = 4'b0001; // x=6, y=23
        pixel_data[23][7] = 4'b0001; // x=7, y=23
        pixel_data[23][8] = 4'b0001; // x=8, y=23
        pixel_data[23][9] = 4'b0001; // x=9, y=23
        pixel_data[23][10] = 4'b0001; // x=10, y=23
        pixel_data[23][11] = 4'b0001; // x=11, y=23
        pixel_data[23][12] = 4'b0001; // x=12, y=23
        pixel_data[23][13] = 4'b0001; // x=13, y=23
        pixel_data[23][14] = 4'b1011; // x=14, y=23
        pixel_data[23][15] = 4'b1011; // x=15, y=23
        pixel_data[23][16] = 4'b0001; // x=16, y=23
        pixel_data[23][17] = 4'b0001; // x=17, y=23
        pixel_data[23][18] = 4'b0001; // x=18, y=23
        pixel_data[23][19] = 4'b0001; // x=19, y=23
        pixel_data[23][20] = 4'b0001; // x=20, y=23
        pixel_data[23][21] = 4'b0001; // x=21, y=23
        pixel_data[23][22] = 4'b0001; // x=22, y=23
        pixel_data[23][23] = 4'b0001; // x=23, y=23
        pixel_data[23][24] = 4'b0001; // x=24, y=23
        pixel_data[23][25] = 4'b0001; // x=25, y=23
        pixel_data[23][26] = 4'b0001; // x=26, y=23
        pixel_data[23][27] = 4'b0001; // x=27, y=23
        pixel_data[23][28] = 4'b0001; // x=28, y=23
        pixel_data[23][29] = 4'b0001; // x=29, y=23
        pixel_data[23][30] = 4'b0001; // x=30, y=23
        pixel_data[23][31] = 4'b1011; // x=31, y=23
        pixel_data[23][32] = 4'b0001; // x=32, y=23
        pixel_data[23][33] = 4'b1101; // x=33, y=23
        pixel_data[23][34] = 4'b1010; // x=34, y=23
        pixel_data[23][35] = 4'b0010; // x=35, y=23
        pixel_data[23][36] = 4'b0010; // x=36, y=23
        pixel_data[23][37] = 4'b0010; // x=37, y=23
        pixel_data[23][38] = 4'b0010; // x=38, y=23
        pixel_data[23][39] = 4'b0010; // x=39, y=23
        pixel_data[23][40] = 4'b0110; // x=40, y=23
        pixel_data[23][41] = 4'b0001; // x=41, y=23
        pixel_data[23][42] = 4'b0001; // x=42, y=23
        pixel_data[23][43] = 4'b0001; // x=43, y=23
        pixel_data[23][44] = 4'b0001; // x=44, y=23
        pixel_data[23][45] = 4'b0001; // x=45, y=23
        pixel_data[23][46] = 4'b0001; // x=46, y=23
        pixel_data[23][47] = 4'b0001; // x=47, y=23
        pixel_data[23][48] = 4'b0001; // x=48, y=23
        pixel_data[23][49] = 4'b0001; // x=49, y=23
        pixel_data[23][50] = 4'b0001; // x=50, y=23
        pixel_data[23][51] = 4'b0001; // x=51, y=23
        pixel_data[23][52] = 4'b0001; // x=52, y=23
        pixel_data[23][53] = 4'b0001; // x=53, y=23
        pixel_data[23][54] = 4'b0001; // x=54, y=23
        pixel_data[23][55] = 4'b0001; // x=55, y=23
        pixel_data[23][56] = 4'b0001; // x=56, y=23
        pixel_data[23][57] = 4'b0001; // x=57, y=23
        pixel_data[23][58] = 4'b0001; // x=58, y=23
        pixel_data[23][59] = 4'b0001; // x=59, y=23
        pixel_data[24][0] = 4'b0001; // x=0, y=24
        pixel_data[24][1] = 4'b0001; // x=1, y=24
        pixel_data[24][2] = 4'b0001; // x=2, y=24
        pixel_data[24][3] = 4'b0001; // x=3, y=24
        pixel_data[24][4] = 4'b0001; // x=4, y=24
        pixel_data[24][5] = 4'b0001; // x=5, y=24
        pixel_data[24][6] = 4'b0001; // x=6, y=24
        pixel_data[24][7] = 4'b0001; // x=7, y=24
        pixel_data[24][8] = 4'b0001; // x=8, y=24
        pixel_data[24][9] = 4'b0001; // x=9, y=24
        pixel_data[24][10] = 4'b0001; // x=10, y=24
        pixel_data[24][11] = 4'b0001; // x=11, y=24
        pixel_data[24][12] = 4'b0001; // x=12, y=24
        pixel_data[24][13] = 4'b0001; // x=13, y=24
        pixel_data[24][14] = 4'b0001; // x=14, y=24
        pixel_data[24][15] = 4'b0001; // x=15, y=24
        pixel_data[24][16] = 4'b0001; // x=16, y=24
        pixel_data[24][17] = 4'b0001; // x=17, y=24
        pixel_data[24][18] = 4'b0001; // x=18, y=24
        pixel_data[24][19] = 4'b0001; // x=19, y=24
        pixel_data[24][20] = 4'b0001; // x=20, y=24
        pixel_data[24][21] = 4'b0001; // x=21, y=24
        pixel_data[24][22] = 4'b0001; // x=22, y=24
        pixel_data[24][23] = 4'b0001; // x=23, y=24
        pixel_data[24][24] = 4'b0001; // x=24, y=24
        pixel_data[24][25] = 4'b0001; // x=25, y=24
        pixel_data[24][26] = 4'b0001; // x=26, y=24
        pixel_data[24][27] = 4'b0001; // x=27, y=24
        pixel_data[24][28] = 4'b0001; // x=28, y=24
        pixel_data[24][29] = 4'b0001; // x=29, y=24
        pixel_data[24][30] = 4'b1011; // x=30, y=24
        pixel_data[24][31] = 4'b0001; // x=31, y=24
        pixel_data[24][32] = 4'b0011; // x=32, y=24
        pixel_data[24][33] = 4'b1010; // x=33, y=24
        pixel_data[24][34] = 4'b0010; // x=34, y=24
        pixel_data[24][35] = 4'b0010; // x=35, y=24
        pixel_data[24][36] = 4'b0010; // x=36, y=24
        pixel_data[24][37] = 4'b0010; // x=37, y=24
        pixel_data[24][38] = 4'b1010; // x=38, y=24
        pixel_data[24][39] = 4'b0101; // x=39, y=24
        pixel_data[24][40] = 4'b0001; // x=40, y=24
        pixel_data[24][41] = 4'b1011; // x=41, y=24
        pixel_data[24][42] = 4'b0001; // x=42, y=24
        pixel_data[24][43] = 4'b0001; // x=43, y=24
        pixel_data[24][44] = 4'b0001; // x=44, y=24
        pixel_data[24][45] = 4'b0001; // x=45, y=24
        pixel_data[24][46] = 4'b0001; // x=46, y=24
        pixel_data[24][47] = 4'b0001; // x=47, y=24
        pixel_data[24][48] = 4'b0001; // x=48, y=24
        pixel_data[24][49] = 4'b0001; // x=49, y=24
        pixel_data[24][50] = 4'b0001; // x=50, y=24
        pixel_data[24][51] = 4'b0001; // x=51, y=24
        pixel_data[24][52] = 4'b0001; // x=52, y=24
        pixel_data[24][53] = 4'b0001; // x=53, y=24
        pixel_data[24][54] = 4'b0001; // x=54, y=24
        pixel_data[24][55] = 4'b0001; // x=55, y=24
        pixel_data[24][56] = 4'b0001; // x=56, y=24
        pixel_data[24][57] = 4'b0001; // x=57, y=24
        pixel_data[24][58] = 4'b0001; // x=58, y=24
        pixel_data[24][59] = 4'b0001; // x=59, y=24
        pixel_data[25][0] = 4'b0001; // x=0, y=25
        pixel_data[25][1] = 4'b0001; // x=1, y=25
        pixel_data[25][2] = 4'b0001; // x=2, y=25
        pixel_data[25][3] = 4'b0001; // x=3, y=25
        pixel_data[25][4] = 4'b0001; // x=4, y=25
        pixel_data[25][5] = 4'b0001; // x=5, y=25
        pixel_data[25][6] = 4'b0001; // x=6, y=25
        pixel_data[25][7] = 4'b0001; // x=7, y=25
        pixel_data[25][8] = 4'b0001; // x=8, y=25
        pixel_data[25][9] = 4'b0001; // x=9, y=25
        pixel_data[25][10] = 4'b0001; // x=10, y=25
        pixel_data[25][11] = 4'b0001; // x=11, y=25
        pixel_data[25][12] = 4'b0001; // x=12, y=25
        pixel_data[25][13] = 4'b0001; // x=13, y=25
        pixel_data[25][14] = 4'b0001; // x=14, y=25
        pixel_data[25][15] = 4'b0001; // x=15, y=25
        pixel_data[25][16] = 4'b0001; // x=16, y=25
        pixel_data[25][17] = 4'b0001; // x=17, y=25
        pixel_data[25][18] = 4'b0001; // x=18, y=25
        pixel_data[25][19] = 4'b0001; // x=19, y=25
        pixel_data[25][20] = 4'b0001; // x=20, y=25
        pixel_data[25][21] = 4'b0001; // x=21, y=25
        pixel_data[25][22] = 4'b0001; // x=22, y=25
        pixel_data[25][23] = 4'b0001; // x=23, y=25
        pixel_data[25][24] = 4'b0001; // x=24, y=25
        pixel_data[25][25] = 4'b0001; // x=25, y=25
        pixel_data[25][26] = 4'b0001; // x=26, y=25
        pixel_data[25][27] = 4'b0001; // x=27, y=25
        pixel_data[25][28] = 4'b0001; // x=28, y=25
        pixel_data[25][29] = 4'b1011; // x=29, y=25
        pixel_data[25][30] = 4'b1011; // x=30, y=25
        pixel_data[25][31] = 4'b1000; // x=31, y=25
        pixel_data[25][32] = 4'b0100; // x=32, y=25
        pixel_data[25][33] = 4'b1010; // x=33, y=25
        pixel_data[25][34] = 4'b0010; // x=34, y=25
        pixel_data[25][35] = 4'b1010; // x=35, y=25
        pixel_data[25][36] = 4'b1010; // x=36, y=25
        pixel_data[25][37] = 4'b1010; // x=37, y=25
        pixel_data[25][38] = 4'b0100; // x=38, y=25
        pixel_data[25][39] = 4'b1110; // x=39, y=25
        pixel_data[25][40] = 4'b1011; // x=40, y=25
        pixel_data[25][41] = 4'b1011; // x=41, y=25
        pixel_data[25][42] = 4'b0001; // x=42, y=25
        pixel_data[25][43] = 4'b0001; // x=43, y=25
        pixel_data[25][44] = 4'b0001; // x=44, y=25
        pixel_data[25][45] = 4'b0001; // x=45, y=25
        pixel_data[25][46] = 4'b0001; // x=46, y=25
        pixel_data[25][47] = 4'b0001; // x=47, y=25
        pixel_data[25][48] = 4'b0001; // x=48, y=25
        pixel_data[25][49] = 4'b0001; // x=49, y=25
        pixel_data[25][50] = 4'b0001; // x=50, y=25
        pixel_data[25][51] = 4'b0001; // x=51, y=25
        pixel_data[25][52] = 4'b0001; // x=52, y=25
        pixel_data[25][53] = 4'b0001; // x=53, y=25
        pixel_data[25][54] = 4'b0001; // x=54, y=25
        pixel_data[25][55] = 4'b0001; // x=55, y=25
        pixel_data[25][56] = 4'b0001; // x=56, y=25
        pixel_data[25][57] = 4'b0001; // x=57, y=25
        pixel_data[25][58] = 4'b0001; // x=58, y=25
        pixel_data[25][59] = 4'b0001; // x=59, y=25
        pixel_data[26][0] = 4'b0001; // x=0, y=26
        pixel_data[26][1] = 4'b0001; // x=1, y=26
        pixel_data[26][2] = 4'b0001; // x=2, y=26
        pixel_data[26][3] = 4'b0001; // x=3, y=26
        pixel_data[26][4] = 4'b0001; // x=4, y=26
        pixel_data[26][5] = 4'b0001; // x=5, y=26
        pixel_data[26][6] = 4'b0001; // x=6, y=26
        pixel_data[26][7] = 4'b0001; // x=7, y=26
        pixel_data[26][8] = 4'b0001; // x=8, y=26
        pixel_data[26][9] = 4'b0001; // x=9, y=26
        pixel_data[26][10] = 4'b0001; // x=10, y=26
        pixel_data[26][11] = 4'b0001; // x=11, y=26
        pixel_data[26][12] = 4'b0001; // x=12, y=26
        pixel_data[26][13] = 4'b0001; // x=13, y=26
        pixel_data[26][14] = 4'b0001; // x=14, y=26
        pixel_data[26][15] = 4'b0001; // x=15, y=26
        pixel_data[26][16] = 4'b0001; // x=16, y=26
        pixel_data[26][17] = 4'b0001; // x=17, y=26
        pixel_data[26][18] = 4'b0001; // x=18, y=26
        pixel_data[26][19] = 4'b0001; // x=19, y=26
        pixel_data[26][20] = 4'b0001; // x=20, y=26
        pixel_data[26][21] = 4'b0001; // x=21, y=26
        pixel_data[26][22] = 4'b0001; // x=22, y=26
        pixel_data[26][23] = 4'b0001; // x=23, y=26
        pixel_data[26][24] = 4'b0001; // x=24, y=26
        pixel_data[26][25] = 4'b0001; // x=25, y=26
        pixel_data[26][26] = 4'b0001; // x=26, y=26
        pixel_data[26][27] = 4'b0001; // x=27, y=26
        pixel_data[26][28] = 4'b0001; // x=28, y=26
        pixel_data[26][29] = 4'b1011; // x=29, y=26
        pixel_data[26][30] = 4'b0001; // x=30, y=26
        pixel_data[26][31] = 4'b0101; // x=31, y=26
        pixel_data[26][32] = 4'b1010; // x=32, y=26
        pixel_data[26][33] = 4'b0010; // x=33, y=26
        pixel_data[26][34] = 4'b1010; // x=34, y=26
        pixel_data[26][35] = 4'b1010; // x=35, y=26
        pixel_data[26][36] = 4'b0010; // x=36, y=26
        pixel_data[26][37] = 4'b1010; // x=37, y=26
        pixel_data[26][38] = 4'b1001; // x=38, y=26
        pixel_data[26][39] = 4'b0001; // x=39, y=26
        pixel_data[26][40] = 4'b1011; // x=40, y=26
        pixel_data[26][41] = 4'b1011; // x=41, y=26
        pixel_data[26][42] = 4'b0001; // x=42, y=26
        pixel_data[26][43] = 4'b0001; // x=43, y=26
        pixel_data[26][44] = 4'b0001; // x=44, y=26
        pixel_data[26][45] = 4'b0001; // x=45, y=26
        pixel_data[26][46] = 4'b0001; // x=46, y=26
        pixel_data[26][47] = 4'b0001; // x=47, y=26
        pixel_data[26][48] = 4'b0001; // x=48, y=26
        pixel_data[26][49] = 4'b0001; // x=49, y=26
        pixel_data[26][50] = 4'b0001; // x=50, y=26
        pixel_data[26][51] = 4'b0001; // x=51, y=26
        pixel_data[26][52] = 4'b0001; // x=52, y=26
        pixel_data[26][53] = 4'b0001; // x=53, y=26
        pixel_data[26][54] = 4'b0001; // x=54, y=26
        pixel_data[26][55] = 4'b0001; // x=55, y=26
        pixel_data[26][56] = 4'b0001; // x=56, y=26
        pixel_data[26][57] = 4'b0001; // x=57, y=26
        pixel_data[26][58] = 4'b0001; // x=58, y=26
        pixel_data[26][59] = 4'b0001; // x=59, y=26
        pixel_data[27][0] = 4'b0001; // x=0, y=27
        pixel_data[27][1] = 4'b0001; // x=1, y=27
        pixel_data[27][2] = 4'b0001; // x=2, y=27
        pixel_data[27][3] = 4'b0001; // x=3, y=27
        pixel_data[27][4] = 4'b0001; // x=4, y=27
        pixel_data[27][5] = 4'b0001; // x=5, y=27
        pixel_data[27][6] = 4'b0001; // x=6, y=27
        pixel_data[27][7] = 4'b0001; // x=7, y=27
        pixel_data[27][8] = 4'b0001; // x=8, y=27
        pixel_data[27][9] = 4'b0001; // x=9, y=27
        pixel_data[27][10] = 4'b0001; // x=10, y=27
        pixel_data[27][11] = 4'b0001; // x=11, y=27
        pixel_data[27][12] = 4'b0001; // x=12, y=27
        pixel_data[27][13] = 4'b0001; // x=13, y=27
        pixel_data[27][14] = 4'b0001; // x=14, y=27
        pixel_data[27][15] = 4'b0001; // x=15, y=27
        pixel_data[27][16] = 4'b0001; // x=16, y=27
        pixel_data[27][17] = 4'b0001; // x=17, y=27
        pixel_data[27][18] = 4'b0001; // x=18, y=27
        pixel_data[27][19] = 4'b0001; // x=19, y=27
        pixel_data[27][20] = 4'b0001; // x=20, y=27
        pixel_data[27][21] = 4'b0001; // x=21, y=27
        pixel_data[27][22] = 4'b0001; // x=22, y=27
        pixel_data[27][23] = 4'b0001; // x=23, y=27
        pixel_data[27][24] = 4'b0001; // x=24, y=27
        pixel_data[27][25] = 4'b0001; // x=25, y=27
        pixel_data[27][26] = 4'b0001; // x=26, y=27
        pixel_data[27][27] = 4'b0001; // x=27, y=27
        pixel_data[27][28] = 4'b1011; // x=28, y=27
        pixel_data[27][29] = 4'b0001; // x=29, y=27
        pixel_data[27][30] = 4'b0110; // x=30, y=27
        pixel_data[27][31] = 4'b0010; // x=31, y=27
        pixel_data[27][32] = 4'b0010; // x=32, y=27
        pixel_data[27][33] = 4'b1010; // x=33, y=27
        pixel_data[27][34] = 4'b1010; // x=34, y=27
        pixel_data[27][35] = 4'b0010; // x=35, y=27
        pixel_data[27][36] = 4'b1010; // x=36, y=27
        pixel_data[27][37] = 4'b0111; // x=37, y=27
        pixel_data[27][38] = 4'b1011; // x=38, y=27
        pixel_data[27][39] = 4'b1011; // x=39, y=27
        pixel_data[27][40] = 4'b1011; // x=40, y=27
        pixel_data[27][41] = 4'b0001; // x=41, y=27
        pixel_data[27][42] = 4'b0001; // x=42, y=27
        pixel_data[27][43] = 4'b0001; // x=43, y=27
        pixel_data[27][44] = 4'b0001; // x=44, y=27
        pixel_data[27][45] = 4'b0001; // x=45, y=27
        pixel_data[27][46] = 4'b0001; // x=46, y=27
        pixel_data[27][47] = 4'b0001; // x=47, y=27
        pixel_data[27][48] = 4'b0001; // x=48, y=27
        pixel_data[27][49] = 4'b0001; // x=49, y=27
        pixel_data[27][50] = 4'b0001; // x=50, y=27
        pixel_data[27][51] = 4'b0001; // x=51, y=27
        pixel_data[27][52] = 4'b0001; // x=52, y=27
        pixel_data[27][53] = 4'b0001; // x=53, y=27
        pixel_data[27][54] = 4'b0001; // x=54, y=27
        pixel_data[27][55] = 4'b0001; // x=55, y=27
        pixel_data[27][56] = 4'b0001; // x=56, y=27
        pixel_data[27][57] = 4'b0001; // x=57, y=27
        pixel_data[27][58] = 4'b0001; // x=58, y=27
        pixel_data[27][59] = 4'b0001; // x=59, y=27
        pixel_data[28][0] = 4'b0001; // x=0, y=28
        pixel_data[28][1] = 4'b0001; // x=1, y=28
        pixel_data[28][2] = 4'b0001; // x=2, y=28
        pixel_data[28][3] = 4'b0001; // x=3, y=28
        pixel_data[28][4] = 4'b0001; // x=4, y=28
        pixel_data[28][5] = 4'b0001; // x=5, y=28
        pixel_data[28][6] = 4'b0001; // x=6, y=28
        pixel_data[28][7] = 4'b0001; // x=7, y=28
        pixel_data[28][8] = 4'b0001; // x=8, y=28
        pixel_data[28][9] = 4'b0001; // x=9, y=28
        pixel_data[28][10] = 4'b0001; // x=10, y=28
        pixel_data[28][11] = 4'b0001; // x=11, y=28
        pixel_data[28][12] = 4'b0001; // x=12, y=28
        pixel_data[28][13] = 4'b0001; // x=13, y=28
        pixel_data[28][14] = 4'b0001; // x=14, y=28
        pixel_data[28][15] = 4'b0001; // x=15, y=28
        pixel_data[28][16] = 4'b0001; // x=16, y=28
        pixel_data[28][17] = 4'b0001; // x=17, y=28
        pixel_data[28][18] = 4'b0001; // x=18, y=28
        pixel_data[28][19] = 4'b0001; // x=19, y=28
        pixel_data[28][20] = 4'b0001; // x=20, y=28
        pixel_data[28][21] = 4'b0001; // x=21, y=28
        pixel_data[28][22] = 4'b0001; // x=22, y=28
        pixel_data[28][23] = 4'b0001; // x=23, y=28
        pixel_data[28][24] = 4'b0001; // x=24, y=28
        pixel_data[28][25] = 4'b0001; // x=25, y=28
        pixel_data[28][26] = 4'b0001; // x=26, y=28
        pixel_data[28][27] = 4'b0001; // x=27, y=28
        pixel_data[28][28] = 4'b1011; // x=28, y=28
        pixel_data[28][29] = 4'b0001; // x=29, y=28
        pixel_data[28][30] = 4'b0111; // x=30, y=28
        pixel_data[28][31] = 4'b1010; // x=31, y=28
        pixel_data[28][32] = 4'b0010; // x=32, y=28
        pixel_data[28][33] = 4'b0010; // x=33, y=28
        pixel_data[28][34] = 4'b0010; // x=34, y=28
        pixel_data[28][35] = 4'b0010; // x=35, y=28
        pixel_data[28][36] = 4'b0010; // x=36, y=28
        pixel_data[28][37] = 4'b1111; // x=37, y=28
        pixel_data[28][38] = 4'b0001; // x=38, y=28
        pixel_data[28][39] = 4'b1011; // x=39, y=28
        pixel_data[28][40] = 4'b0001; // x=40, y=28
        pixel_data[28][41] = 4'b0001; // x=41, y=28
        pixel_data[28][42] = 4'b0001; // x=42, y=28
        pixel_data[28][43] = 4'b0001; // x=43, y=28
        pixel_data[28][44] = 4'b0001; // x=44, y=28
        pixel_data[28][45] = 4'b0001; // x=45, y=28
        pixel_data[28][46] = 4'b0001; // x=46, y=28
        pixel_data[28][47] = 4'b0001; // x=47, y=28
        pixel_data[28][48] = 4'b0001; // x=48, y=28
        pixel_data[28][49] = 4'b0001; // x=49, y=28
        pixel_data[28][50] = 4'b0001; // x=50, y=28
        pixel_data[28][51] = 4'b0001; // x=51, y=28
        pixel_data[28][52] = 4'b0001; // x=52, y=28
        pixel_data[28][53] = 4'b0001; // x=53, y=28
        pixel_data[28][54] = 4'b0001; // x=54, y=28
        pixel_data[28][55] = 4'b0001; // x=55, y=28
        pixel_data[28][56] = 4'b0001; // x=56, y=28
        pixel_data[28][57] = 4'b0001; // x=57, y=28
        pixel_data[28][58] = 4'b0001; // x=58, y=28
        pixel_data[28][59] = 4'b0001; // x=59, y=28
        pixel_data[29][0] = 4'b0001; // x=0, y=29
        pixel_data[29][1] = 4'b0001; // x=1, y=29
        pixel_data[29][2] = 4'b0001; // x=2, y=29
        pixel_data[29][3] = 4'b0001; // x=3, y=29
        pixel_data[29][4] = 4'b0001; // x=4, y=29
        pixel_data[29][5] = 4'b0001; // x=5, y=29
        pixel_data[29][6] = 4'b0001; // x=6, y=29
        pixel_data[29][7] = 4'b0001; // x=7, y=29
        pixel_data[29][8] = 4'b0001; // x=8, y=29
        pixel_data[29][9] = 4'b0001; // x=9, y=29
        pixel_data[29][10] = 4'b0001; // x=10, y=29
        pixel_data[29][11] = 4'b0001; // x=11, y=29
        pixel_data[29][12] = 4'b0001; // x=12, y=29
        pixel_data[29][13] = 4'b0001; // x=13, y=29
        pixel_data[29][14] = 4'b0001; // x=14, y=29
        pixel_data[29][15] = 4'b0001; // x=15, y=29
        pixel_data[29][16] = 4'b0001; // x=16, y=29
        pixel_data[29][17] = 4'b0001; // x=17, y=29
        pixel_data[29][18] = 4'b0001; // x=18, y=29
        pixel_data[29][19] = 4'b0001; // x=19, y=29
        pixel_data[29][20] = 4'b0001; // x=20, y=29
        pixel_data[29][21] = 4'b0001; // x=21, y=29
        pixel_data[29][22] = 4'b0001; // x=22, y=29
        pixel_data[29][23] = 4'b0001; // x=23, y=29
        pixel_data[29][24] = 4'b0001; // x=24, y=29
        pixel_data[29][25] = 4'b0001; // x=25, y=29
        pixel_data[29][26] = 4'b0001; // x=26, y=29
        pixel_data[29][27] = 4'b0001; // x=27, y=29
        pixel_data[29][28] = 4'b0001; // x=28, y=29
        pixel_data[29][29] = 4'b0011; // x=29, y=29
        pixel_data[29][30] = 4'b1010; // x=30, y=29
        pixel_data[29][31] = 4'b0010; // x=31, y=29
        pixel_data[29][32] = 4'b0010; // x=32, y=29
        pixel_data[29][33] = 4'b0010; // x=33, y=29
        pixel_data[29][34] = 4'b0010; // x=34, y=29
        pixel_data[29][35] = 4'b1010; // x=35, y=29
        pixel_data[29][36] = 4'b1101; // x=36, y=29
        pixel_data[29][37] = 4'b0001; // x=37, y=29
        pixel_data[29][38] = 4'b0001; // x=38, y=29
        pixel_data[29][39] = 4'b0001; // x=39, y=29
        pixel_data[29][40] = 4'b0001; // x=40, y=29
        pixel_data[29][41] = 4'b0001; // x=41, y=29
        pixel_data[29][42] = 4'b0001; // x=42, y=29
        pixel_data[29][43] = 4'b0001; // x=43, y=29
        pixel_data[29][44] = 4'b0001; // x=44, y=29
        pixel_data[29][45] = 4'b0001; // x=45, y=29
        pixel_data[29][46] = 4'b0001; // x=46, y=29
        pixel_data[29][47] = 4'b0001; // x=47, y=29
        pixel_data[29][48] = 4'b0001; // x=48, y=29
        pixel_data[29][49] = 4'b0001; // x=49, y=29
        pixel_data[29][50] = 4'b0001; // x=50, y=29
        pixel_data[29][51] = 4'b0001; // x=51, y=29
        pixel_data[29][52] = 4'b0001; // x=52, y=29
        pixel_data[29][53] = 4'b0001; // x=53, y=29
        pixel_data[29][54] = 4'b0001; // x=54, y=29
        pixel_data[29][55] = 4'b0001; // x=55, y=29
        pixel_data[29][56] = 4'b0001; // x=56, y=29
        pixel_data[29][57] = 4'b0001; // x=57, y=29
        pixel_data[29][58] = 4'b0001; // x=58, y=29
        pixel_data[29][59] = 4'b0001; // x=59, y=29
        pixel_data[30][0] = 4'b0001; // x=0, y=30
        pixel_data[30][1] = 4'b0001; // x=1, y=30
        pixel_data[30][2] = 4'b0001; // x=2, y=30
        pixel_data[30][3] = 4'b0001; // x=3, y=30
        pixel_data[30][4] = 4'b0001; // x=4, y=30
        pixel_data[30][5] = 4'b0001; // x=5, y=30
        pixel_data[30][6] = 4'b0001; // x=6, y=30
        pixel_data[30][7] = 4'b0001; // x=7, y=30
        pixel_data[30][8] = 4'b0001; // x=8, y=30
        pixel_data[30][9] = 4'b0001; // x=9, y=30
        pixel_data[30][10] = 4'b0001; // x=10, y=30
        pixel_data[30][11] = 4'b0001; // x=11, y=30
        pixel_data[30][12] = 4'b0001; // x=12, y=30
        pixel_data[30][13] = 4'b0001; // x=13, y=30
        pixel_data[30][14] = 4'b0001; // x=14, y=30
        pixel_data[30][15] = 4'b0001; // x=15, y=30
        pixel_data[30][16] = 4'b0001; // x=16, y=30
        pixel_data[30][17] = 4'b0001; // x=17, y=30
        pixel_data[30][18] = 4'b0001; // x=18, y=30
        pixel_data[30][19] = 4'b0001; // x=19, y=30
        pixel_data[30][20] = 4'b0001; // x=20, y=30
        pixel_data[30][21] = 4'b0001; // x=21, y=30
        pixel_data[30][22] = 4'b0001; // x=22, y=30
        pixel_data[30][23] = 4'b0001; // x=23, y=30
        pixel_data[30][24] = 4'b0001; // x=24, y=30
        pixel_data[30][25] = 4'b0001; // x=25, y=30
        pixel_data[30][26] = 4'b0001; // x=26, y=30
        pixel_data[30][27] = 4'b0001; // x=27, y=30
        pixel_data[30][28] = 4'b1000; // x=28, y=30
        pixel_data[30][29] = 4'b0100; // x=29, y=30
        pixel_data[30][30] = 4'b1010; // x=30, y=30
        pixel_data[30][31] = 4'b0010; // x=31, y=30
        pixel_data[30][32] = 4'b0010; // x=32, y=30
        pixel_data[30][33] = 4'b0010; // x=33, y=30
        pixel_data[30][34] = 4'b1010; // x=34, y=30
        pixel_data[30][35] = 4'b0100; // x=35, y=30
        pixel_data[30][36] = 4'b1110; // x=36, y=30
        pixel_data[30][37] = 4'b0001; // x=37, y=30
        pixel_data[30][38] = 4'b0001; // x=38, y=30
        pixel_data[30][39] = 4'b0001; // x=39, y=30
        pixel_data[30][40] = 4'b0001; // x=40, y=30
        pixel_data[30][41] = 4'b0001; // x=41, y=30
        pixel_data[30][42] = 4'b0001; // x=42, y=30
        pixel_data[30][43] = 4'b0001; // x=43, y=30
        pixel_data[30][44] = 4'b0001; // x=44, y=30
        pixel_data[30][45] = 4'b0001; // x=45, y=30
        pixel_data[30][46] = 4'b0001; // x=46, y=30
        pixel_data[30][47] = 4'b0001; // x=47, y=30
        pixel_data[30][48] = 4'b0001; // x=48, y=30
        pixel_data[30][49] = 4'b0001; // x=49, y=30
        pixel_data[30][50] = 4'b0001; // x=50, y=30
        pixel_data[30][51] = 4'b0001; // x=51, y=30
        pixel_data[30][52] = 4'b0001; // x=52, y=30
        pixel_data[30][53] = 4'b0001; // x=53, y=30
        pixel_data[30][54] = 4'b0001; // x=54, y=30
        pixel_data[30][55] = 4'b0001; // x=55, y=30
        pixel_data[30][56] = 4'b0001; // x=56, y=30
        pixel_data[30][57] = 4'b0001; // x=57, y=30
        pixel_data[30][58] = 4'b0001; // x=58, y=30
        pixel_data[30][59] = 4'b0001; // x=59, y=30
        pixel_data[31][0] = 4'b0001; // x=0, y=31
        pixel_data[31][1] = 4'b0001; // x=1, y=31
        pixel_data[31][2] = 4'b0001; // x=2, y=31
        pixel_data[31][3] = 4'b0001; // x=3, y=31
        pixel_data[31][4] = 4'b0001; // x=4, y=31
        pixel_data[31][5] = 4'b0001; // x=5, y=31
        pixel_data[31][6] = 4'b0001; // x=6, y=31
        pixel_data[31][7] = 4'b0001; // x=7, y=31
        pixel_data[31][8] = 4'b0001; // x=8, y=31
        pixel_data[31][9] = 4'b0001; // x=9, y=31
        pixel_data[31][10] = 4'b0001; // x=10, y=31
        pixel_data[31][11] = 4'b0001; // x=11, y=31
        pixel_data[31][12] = 4'b0001; // x=12, y=31
        pixel_data[31][13] = 4'b0001; // x=13, y=31
        pixel_data[31][14] = 4'b0001; // x=14, y=31
        pixel_data[31][15] = 4'b0001; // x=15, y=31
        pixel_data[31][16] = 4'b0001; // x=16, y=31
        pixel_data[31][17] = 4'b0001; // x=17, y=31
        pixel_data[31][18] = 4'b0001; // x=18, y=31
        pixel_data[31][19] = 4'b0001; // x=19, y=31
        pixel_data[31][20] = 4'b0001; // x=20, y=31
        pixel_data[31][21] = 4'b0001; // x=21, y=31
        pixel_data[31][22] = 4'b0001; // x=22, y=31
        pixel_data[31][23] = 4'b0001; // x=23, y=31
        pixel_data[31][24] = 4'b0001; // x=24, y=31
        pixel_data[31][25] = 4'b0001; // x=25, y=31
        pixel_data[31][26] = 4'b1011; // x=26, y=31
        pixel_data[31][27] = 4'b0001; // x=27, y=31
        pixel_data[31][28] = 4'b0101; // x=28, y=31
        pixel_data[31][29] = 4'b1010; // x=29, y=31
        pixel_data[31][30] = 4'b0010; // x=30, y=31
        pixel_data[31][31] = 4'b1010; // x=31, y=31
        pixel_data[31][32] = 4'b1010; // x=32, y=31
        pixel_data[31][33] = 4'b0010; // x=33, y=31
        pixel_data[31][34] = 4'b1010; // x=34, y=31
        pixel_data[31][35] = 4'b1100; // x=35, y=31
        pixel_data[31][36] = 4'b0001; // x=36, y=31
        pixel_data[31][37] = 4'b1011; // x=37, y=31
        pixel_data[31][38] = 4'b0001; // x=38, y=31
        pixel_data[31][39] = 4'b0001; // x=39, y=31
        pixel_data[31][40] = 4'b0001; // x=40, y=31
        pixel_data[31][41] = 4'b0001; // x=41, y=31
        pixel_data[31][42] = 4'b0001; // x=42, y=31
        pixel_data[31][43] = 4'b0001; // x=43, y=31
        pixel_data[31][44] = 4'b0001; // x=44, y=31
        pixel_data[31][45] = 4'b0001; // x=45, y=31
        pixel_data[31][46] = 4'b0001; // x=46, y=31
        pixel_data[31][47] = 4'b0001; // x=47, y=31
        pixel_data[31][48] = 4'b0001; // x=48, y=31
        pixel_data[31][49] = 4'b0001; // x=49, y=31
        pixel_data[31][50] = 4'b0001; // x=50, y=31
        pixel_data[31][51] = 4'b0001; // x=51, y=31
        pixel_data[31][52] = 4'b0001; // x=52, y=31
        pixel_data[31][53] = 4'b0001; // x=53, y=31
        pixel_data[31][54] = 4'b0001; // x=54, y=31
        pixel_data[31][55] = 4'b0001; // x=55, y=31
        pixel_data[31][56] = 4'b0001; // x=56, y=31
        pixel_data[31][57] = 4'b0001; // x=57, y=31
        pixel_data[31][58] = 4'b0001; // x=58, y=31
        pixel_data[31][59] = 4'b0001; // x=59, y=31
        pixel_data[32][0] = 4'b0001; // x=0, y=32
        pixel_data[32][1] = 4'b0001; // x=1, y=32
        pixel_data[32][2] = 4'b0001; // x=2, y=32
        pixel_data[32][3] = 4'b0001; // x=3, y=32
        pixel_data[32][4] = 4'b0001; // x=4, y=32
        pixel_data[32][5] = 4'b0001; // x=5, y=32
        pixel_data[32][6] = 4'b0001; // x=6, y=32
        pixel_data[32][7] = 4'b0001; // x=7, y=32
        pixel_data[32][8] = 4'b0001; // x=8, y=32
        pixel_data[32][9] = 4'b0001; // x=9, y=32
        pixel_data[32][10] = 4'b0001; // x=10, y=32
        pixel_data[32][11] = 4'b0001; // x=11, y=32
        pixel_data[32][12] = 4'b0001; // x=12, y=32
        pixel_data[32][13] = 4'b0001; // x=13, y=32
        pixel_data[32][14] = 4'b0001; // x=14, y=32
        pixel_data[32][15] = 4'b0001; // x=15, y=32
        pixel_data[32][16] = 4'b0001; // x=16, y=32
        pixel_data[32][17] = 4'b0001; // x=17, y=32
        pixel_data[32][18] = 4'b0001; // x=18, y=32
        pixel_data[32][19] = 4'b0001; // x=19, y=32
        pixel_data[32][20] = 4'b0001; // x=20, y=32
        pixel_data[32][21] = 4'b0001; // x=21, y=32
        pixel_data[32][22] = 4'b0001; // x=22, y=32
        pixel_data[32][23] = 4'b0001; // x=23, y=32
        pixel_data[32][24] = 4'b0001; // x=24, y=32
        pixel_data[32][25] = 4'b1011; // x=25, y=32
        pixel_data[32][26] = 4'b0001; // x=26, y=32
        pixel_data[32][27] = 4'b0110; // x=27, y=32
        pixel_data[32][28] = 4'b0010; // x=28, y=32
        pixel_data[32][29] = 4'b0010; // x=29, y=32
        pixel_data[32][30] = 4'b1010; // x=30, y=32
        pixel_data[32][31] = 4'b1010; // x=31, y=32
        pixel_data[32][32] = 4'b1010; // x=32, y=32
        pixel_data[32][33] = 4'b1010; // x=33, y=32
        pixel_data[32][34] = 4'b0000; // x=34, y=32
        pixel_data[32][35] = 4'b1000; // x=35, y=32
        pixel_data[32][36] = 4'b1011; // x=36, y=32
        pixel_data[32][37] = 4'b0001; // x=37, y=32
        pixel_data[32][38] = 4'b0001; // x=38, y=32
        pixel_data[32][39] = 4'b0001; // x=39, y=32
        pixel_data[32][40] = 4'b0001; // x=40, y=32
        pixel_data[32][41] = 4'b0001; // x=41, y=32
        pixel_data[32][42] = 4'b0001; // x=42, y=32
        pixel_data[32][43] = 4'b0001; // x=43, y=32
        pixel_data[32][44] = 4'b0001; // x=44, y=32
        pixel_data[32][45] = 4'b0001; // x=45, y=32
        pixel_data[32][46] = 4'b0001; // x=46, y=32
        pixel_data[32][47] = 4'b0001; // x=47, y=32
        pixel_data[32][48] = 4'b0001; // x=48, y=32
        pixel_data[32][49] = 4'b0001; // x=49, y=32
        pixel_data[32][50] = 4'b0001; // x=50, y=32
        pixel_data[32][51] = 4'b0001; // x=51, y=32
        pixel_data[32][52] = 4'b0001; // x=52, y=32
        pixel_data[32][53] = 4'b0001; // x=53, y=32
        pixel_data[32][54] = 4'b0001; // x=54, y=32
        pixel_data[32][55] = 4'b0001; // x=55, y=32
        pixel_data[32][56] = 4'b0001; // x=56, y=32
        pixel_data[32][57] = 4'b0001; // x=57, y=32
        pixel_data[32][58] = 4'b0001; // x=58, y=32
        pixel_data[32][59] = 4'b0001; // x=59, y=32
        pixel_data[33][0] = 4'b0001; // x=0, y=33
        pixel_data[33][1] = 4'b0001; // x=1, y=33
        pixel_data[33][2] = 4'b0001; // x=2, y=33
        pixel_data[33][3] = 4'b0001; // x=3, y=33
        pixel_data[33][4] = 4'b0001; // x=4, y=33
        pixel_data[33][5] = 4'b0001; // x=5, y=33
        pixel_data[33][6] = 4'b0001; // x=6, y=33
        pixel_data[33][7] = 4'b0001; // x=7, y=33
        pixel_data[33][8] = 4'b0001; // x=8, y=33
        pixel_data[33][9] = 4'b0001; // x=9, y=33
        pixel_data[33][10] = 4'b0001; // x=10, y=33
        pixel_data[33][11] = 4'b0001; // x=11, y=33
        pixel_data[33][12] = 4'b0001; // x=12, y=33
        pixel_data[33][13] = 4'b0001; // x=13, y=33
        pixel_data[33][14] = 4'b0001; // x=14, y=33
        pixel_data[33][15] = 4'b0001; // x=15, y=33
        pixel_data[33][16] = 4'b0001; // x=16, y=33
        pixel_data[33][17] = 4'b0001; // x=17, y=33
        pixel_data[33][18] = 4'b0001; // x=18, y=33
        pixel_data[33][19] = 4'b0001; // x=19, y=33
        pixel_data[33][20] = 4'b0001; // x=20, y=33
        pixel_data[33][21] = 4'b0001; // x=21, y=33
        pixel_data[33][22] = 4'b0001; // x=22, y=33
        pixel_data[33][23] = 4'b0001; // x=23, y=33
        pixel_data[33][24] = 4'b1011; // x=24, y=33
        pixel_data[33][25] = 4'b1011; // x=25, y=33
        pixel_data[33][26] = 4'b1011; // x=26, y=33
        pixel_data[33][27] = 4'b0111; // x=27, y=33
        pixel_data[33][28] = 4'b1010; // x=28, y=33
        pixel_data[33][29] = 4'b0010; // x=29, y=33
        pixel_data[33][30] = 4'b1010; // x=30, y=33
        pixel_data[33][31] = 4'b1010; // x=31, y=33
        pixel_data[33][32] = 4'b0010; // x=32, y=33
        pixel_data[33][33] = 4'b1010; // x=33, y=33
        pixel_data[33][34] = 4'b0011; // x=34, y=33
        pixel_data[33][35] = 4'b0001; // x=35, y=33
        pixel_data[33][36] = 4'b1011; // x=36, y=33
        pixel_data[33][37] = 4'b0001; // x=37, y=33
        pixel_data[33][38] = 4'b0001; // x=38, y=33
        pixel_data[33][39] = 4'b0001; // x=39, y=33
        pixel_data[33][40] = 4'b0001; // x=40, y=33
        pixel_data[33][41] = 4'b0001; // x=41, y=33
        pixel_data[33][42] = 4'b0001; // x=42, y=33
        pixel_data[33][43] = 4'b0001; // x=43, y=33
        pixel_data[33][44] = 4'b0001; // x=44, y=33
        pixel_data[33][45] = 4'b0001; // x=45, y=33
        pixel_data[33][46] = 4'b0001; // x=46, y=33
        pixel_data[33][47] = 4'b0001; // x=47, y=33
        pixel_data[33][48] = 4'b0001; // x=48, y=33
        pixel_data[33][49] = 4'b0001; // x=49, y=33
        pixel_data[33][50] = 4'b0001; // x=50, y=33
        pixel_data[33][51] = 4'b0001; // x=51, y=33
        pixel_data[33][52] = 4'b0001; // x=52, y=33
        pixel_data[33][53] = 4'b0001; // x=53, y=33
        pixel_data[33][54] = 4'b0001; // x=54, y=33
        pixel_data[33][55] = 4'b0001; // x=55, y=33
        pixel_data[33][56] = 4'b0001; // x=56, y=33
        pixel_data[33][57] = 4'b0001; // x=57, y=33
        pixel_data[33][58] = 4'b0001; // x=58, y=33
        pixel_data[33][59] = 4'b0001; // x=59, y=33
        pixel_data[34][0] = 4'b0001; // x=0, y=34
        pixel_data[34][1] = 4'b0001; // x=1, y=34
        pixel_data[34][2] = 4'b0001; // x=2, y=34
        pixel_data[34][3] = 4'b0001; // x=3, y=34
        pixel_data[34][4] = 4'b0001; // x=4, y=34
        pixel_data[34][5] = 4'b0001; // x=5, y=34
        pixel_data[34][6] = 4'b0001; // x=6, y=34
        pixel_data[34][7] = 4'b0001; // x=7, y=34
        pixel_data[34][8] = 4'b0001; // x=8, y=34
        pixel_data[34][9] = 4'b0001; // x=9, y=34
        pixel_data[34][10] = 4'b0001; // x=10, y=34
        pixel_data[34][11] = 4'b0001; // x=11, y=34
        pixel_data[34][12] = 4'b0001; // x=12, y=34
        pixel_data[34][13] = 4'b0001; // x=13, y=34
        pixel_data[34][14] = 4'b0001; // x=14, y=34
        pixel_data[34][15] = 4'b0001; // x=15, y=34
        pixel_data[34][16] = 4'b0001; // x=16, y=34
        pixel_data[34][17] = 4'b0001; // x=17, y=34
        pixel_data[34][18] = 4'b0001; // x=18, y=34
        pixel_data[34][19] = 4'b0001; // x=19, y=34
        pixel_data[34][20] = 4'b0001; // x=20, y=34
        pixel_data[34][21] = 4'b0001; // x=21, y=34
        pixel_data[34][22] = 4'b0001; // x=22, y=34
        pixel_data[34][23] = 4'b0001; // x=23, y=34
        pixel_data[34][24] = 4'b1011; // x=24, y=34
        pixel_data[34][25] = 4'b0001; // x=25, y=34
        pixel_data[34][26] = 4'b1001; // x=26, y=34
        pixel_data[34][27] = 4'b1010; // x=27, y=34
        pixel_data[34][28] = 4'b1010; // x=28, y=34
        pixel_data[34][29] = 4'b1010; // x=29, y=34
        pixel_data[34][30] = 4'b1010; // x=30, y=34
        pixel_data[34][31] = 4'b0010; // x=31, y=34
        pixel_data[34][32] = 4'b1010; // x=32, y=34
        pixel_data[34][33] = 4'b1101; // x=33, y=34
        pixel_data[34][34] = 4'b0001; // x=34, y=34
        pixel_data[34][35] = 4'b1011; // x=35, y=34
        pixel_data[34][36] = 4'b1011; // x=36, y=34
        pixel_data[34][37] = 4'b1011; // x=37, y=34
        pixel_data[34][38] = 4'b0001; // x=38, y=34
        pixel_data[34][39] = 4'b0001; // x=39, y=34
        pixel_data[34][40] = 4'b0001; // x=40, y=34
        pixel_data[34][41] = 4'b0001; // x=41, y=34
        pixel_data[34][42] = 4'b0001; // x=42, y=34
        pixel_data[34][43] = 4'b0001; // x=43, y=34
        pixel_data[34][44] = 4'b0001; // x=44, y=34
        pixel_data[34][45] = 4'b0001; // x=45, y=34
        pixel_data[34][46] = 4'b0001; // x=46, y=34
        pixel_data[34][47] = 4'b0001; // x=47, y=34
        pixel_data[34][48] = 4'b0001; // x=48, y=34
        pixel_data[34][49] = 4'b0001; // x=49, y=34
        pixel_data[34][50] = 4'b0001; // x=50, y=34
        pixel_data[34][51] = 4'b0001; // x=51, y=34
        pixel_data[34][52] = 4'b0001; // x=52, y=34
        pixel_data[34][53] = 4'b0001; // x=53, y=34
        pixel_data[34][54] = 4'b0001; // x=54, y=34
        pixel_data[34][55] = 4'b0001; // x=55, y=34
        pixel_data[34][56] = 4'b0001; // x=56, y=34
        pixel_data[34][57] = 4'b0001; // x=57, y=34
        pixel_data[34][58] = 4'b0001; // x=58, y=34
        pixel_data[34][59] = 4'b0001; // x=59, y=34
        pixel_data[35][0] = 4'b0001; // x=0, y=35
        pixel_data[35][1] = 4'b0001; // x=1, y=35
        pixel_data[35][2] = 4'b0001; // x=2, y=35
        pixel_data[35][3] = 4'b0001; // x=3, y=35
        pixel_data[35][4] = 4'b0001; // x=4, y=35
        pixel_data[35][5] = 4'b0001; // x=5, y=35
        pixel_data[35][6] = 4'b0001; // x=6, y=35
        pixel_data[35][7] = 4'b0001; // x=7, y=35
        pixel_data[35][8] = 4'b0001; // x=8, y=35
        pixel_data[35][9] = 4'b0001; // x=9, y=35
        pixel_data[35][10] = 4'b0001; // x=10, y=35
        pixel_data[35][11] = 4'b0001; // x=11, y=35
        pixel_data[35][12] = 4'b0001; // x=12, y=35
        pixel_data[35][13] = 4'b0001; // x=13, y=35
        pixel_data[35][14] = 4'b0001; // x=14, y=35
        pixel_data[35][15] = 4'b0001; // x=15, y=35
        pixel_data[35][16] = 4'b0001; // x=16, y=35
        pixel_data[35][17] = 4'b0001; // x=17, y=35
        pixel_data[35][18] = 4'b0001; // x=18, y=35
        pixel_data[35][19] = 4'b0001; // x=19, y=35
        pixel_data[35][20] = 4'b0001; // x=20, y=35
        pixel_data[35][21] = 4'b0001; // x=21, y=35
        pixel_data[35][22] = 4'b0001; // x=22, y=35
        pixel_data[35][23] = 4'b0001; // x=23, y=35
        pixel_data[35][24] = 4'b0001; // x=24, y=35
        pixel_data[35][25] = 4'b1110; // x=25, y=35
        pixel_data[35][26] = 4'b0100; // x=26, y=35
        pixel_data[35][27] = 4'b1010; // x=27, y=35
        pixel_data[35][28] = 4'b0010; // x=28, y=35
        pixel_data[35][29] = 4'b1010; // x=29, y=35
        pixel_data[35][30] = 4'b1010; // x=30, y=35
        pixel_data[35][31] = 4'b1010; // x=31, y=35
        pixel_data[35][32] = 4'b0010; // x=32, y=35
        pixel_data[35][33] = 4'b0110; // x=33, y=35
        pixel_data[35][34] = 4'b0001; // x=34, y=35
        pixel_data[35][35] = 4'b1011; // x=35, y=35
        pixel_data[35][36] = 4'b0001; // x=36, y=35
        pixel_data[35][37] = 4'b0001; // x=37, y=35
        pixel_data[35][38] = 4'b0001; // x=38, y=35
        pixel_data[35][39] = 4'b0001; // x=39, y=35
        pixel_data[35][40] = 4'b0001; // x=40, y=35
        pixel_data[35][41] = 4'b0001; // x=41, y=35
        pixel_data[35][42] = 4'b0001; // x=42, y=35
        pixel_data[35][43] = 4'b0001; // x=43, y=35
        pixel_data[35][44] = 4'b0001; // x=44, y=35
        pixel_data[35][45] = 4'b0001; // x=45, y=35
        pixel_data[35][46] = 4'b0001; // x=46, y=35
        pixel_data[35][47] = 4'b0001; // x=47, y=35
        pixel_data[35][48] = 4'b0001; // x=48, y=35
        pixel_data[35][49] = 4'b0001; // x=49, y=35
        pixel_data[35][50] = 4'b0001; // x=50, y=35
        pixel_data[35][51] = 4'b0001; // x=51, y=35
        pixel_data[35][52] = 4'b0001; // x=52, y=35
        pixel_data[35][53] = 4'b0001; // x=53, y=35
        pixel_data[35][54] = 4'b0001; // x=54, y=35
        pixel_data[35][55] = 4'b0001; // x=55, y=35
        pixel_data[35][56] = 4'b0001; // x=56, y=35
        pixel_data[35][57] = 4'b0001; // x=57, y=35
        pixel_data[35][58] = 4'b0001; // x=58, y=35
        pixel_data[35][59] = 4'b0001; // x=59, y=35
        pixel_data[36][0] = 4'b0001; // x=0, y=36
        pixel_data[36][1] = 4'b0001; // x=1, y=36
        pixel_data[36][2] = 4'b0001; // x=2, y=36
        pixel_data[36][3] = 4'b0001; // x=3, y=36
        pixel_data[36][4] = 4'b0001; // x=4, y=36
        pixel_data[36][5] = 4'b0001; // x=5, y=36
        pixel_data[36][6] = 4'b0001; // x=6, y=36
        pixel_data[36][7] = 4'b0001; // x=7, y=36
        pixel_data[36][8] = 4'b0001; // x=8, y=36
        pixel_data[36][9] = 4'b0001; // x=9, y=36
        pixel_data[36][10] = 4'b0001; // x=10, y=36
        pixel_data[36][11] = 4'b0001; // x=11, y=36
        pixel_data[36][12] = 4'b0001; // x=12, y=36
        pixel_data[36][13] = 4'b0001; // x=13, y=36
        pixel_data[36][14] = 4'b0001; // x=14, y=36
        pixel_data[36][15] = 4'b0001; // x=15, y=36
        pixel_data[36][16] = 4'b0001; // x=16, y=36
        pixel_data[36][17] = 4'b0001; // x=17, y=36
        pixel_data[36][18] = 4'b0001; // x=18, y=36
        pixel_data[36][19] = 4'b0001; // x=19, y=36
        pixel_data[36][20] = 4'b0001; // x=20, y=36
        pixel_data[36][21] = 4'b0001; // x=21, y=36
        pixel_data[36][22] = 4'b0001; // x=22, y=36
        pixel_data[36][23] = 4'b1011; // x=23, y=36
        pixel_data[36][24] = 4'b0001; // x=24, y=36
        pixel_data[36][25] = 4'b0101; // x=25, y=36
        pixel_data[36][26] = 4'b1010; // x=26, y=36
        pixel_data[36][27] = 4'b0010; // x=27, y=36
        pixel_data[36][28] = 4'b0010; // x=28, y=36
        pixel_data[36][29] = 4'b1010; // x=29, y=36
        pixel_data[36][30] = 4'b0010; // x=30, y=36
        pixel_data[36][31] = 4'b1010; // x=31, y=36
        pixel_data[36][32] = 4'b0101; // x=32, y=36
        pixel_data[36][33] = 4'b0001; // x=33, y=36
        pixel_data[36][34] = 4'b1011; // x=34, y=36
        pixel_data[36][35] = 4'b0001; // x=35, y=36
        pixel_data[36][36] = 4'b0001; // x=36, y=36
        pixel_data[36][37] = 4'b0001; // x=37, y=36
        pixel_data[36][38] = 4'b0001; // x=38, y=36
        pixel_data[36][39] = 4'b0001; // x=39, y=36
        pixel_data[36][40] = 4'b0001; // x=40, y=36
        pixel_data[36][41] = 4'b0001; // x=41, y=36
        pixel_data[36][42] = 4'b0001; // x=42, y=36
        pixel_data[36][43] = 4'b0001; // x=43, y=36
        pixel_data[36][44] = 4'b0001; // x=44, y=36
        pixel_data[36][45] = 4'b0001; // x=45, y=36
        pixel_data[36][46] = 4'b0001; // x=46, y=36
        pixel_data[36][47] = 4'b0001; // x=47, y=36
        pixel_data[36][48] = 4'b0001; // x=48, y=36
        pixel_data[36][49] = 4'b0001; // x=49, y=36
        pixel_data[36][50] = 4'b0001; // x=50, y=36
        pixel_data[36][51] = 4'b0001; // x=51, y=36
        pixel_data[36][52] = 4'b0001; // x=52, y=36
        pixel_data[36][53] = 4'b0001; // x=53, y=36
        pixel_data[36][54] = 4'b0001; // x=54, y=36
        pixel_data[36][55] = 4'b0001; // x=55, y=36
        pixel_data[36][56] = 4'b0001; // x=56, y=36
        pixel_data[36][57] = 4'b0001; // x=57, y=36
        pixel_data[36][58] = 4'b0001; // x=58, y=36
        pixel_data[36][59] = 4'b0001; // x=59, y=36
        pixel_data[37][0] = 4'b0001; // x=0, y=37
        pixel_data[37][1] = 4'b0001; // x=1, y=37
        pixel_data[37][2] = 4'b0001; // x=2, y=37
        pixel_data[37][3] = 4'b0001; // x=3, y=37
        pixel_data[37][4] = 4'b0001; // x=4, y=37
        pixel_data[37][5] = 4'b0001; // x=5, y=37
        pixel_data[37][6] = 4'b0001; // x=6, y=37
        pixel_data[37][7] = 4'b0001; // x=7, y=37
        pixel_data[37][8] = 4'b0001; // x=8, y=37
        pixel_data[37][9] = 4'b0001; // x=9, y=37
        pixel_data[37][10] = 4'b0001; // x=10, y=37
        pixel_data[37][11] = 4'b0001; // x=11, y=37
        pixel_data[37][12] = 4'b0001; // x=12, y=37
        pixel_data[37][13] = 4'b0001; // x=13, y=37
        pixel_data[37][14] = 4'b0001; // x=14, y=37
        pixel_data[37][15] = 4'b0001; // x=15, y=37
        pixel_data[37][16] = 4'b0001; // x=16, y=37
        pixel_data[37][17] = 4'b0001; // x=17, y=37
        pixel_data[37][18] = 4'b0001; // x=18, y=37
        pixel_data[37][19] = 4'b0001; // x=19, y=37
        pixel_data[37][20] = 4'b0001; // x=20, y=37
        pixel_data[37][21] = 4'b0001; // x=21, y=37
        pixel_data[37][22] = 4'b0001; // x=22, y=37
        pixel_data[37][23] = 4'b0001; // x=23, y=37
        pixel_data[37][24] = 4'b0110; // x=24, y=37
        pixel_data[37][25] = 4'b0010; // x=25, y=37
        pixel_data[37][26] = 4'b1010; // x=26, y=37
        pixel_data[37][27] = 4'b1010; // x=27, y=37
        pixel_data[37][28] = 4'b0010; // x=28, y=37
        pixel_data[37][29] = 4'b0010; // x=29, y=37
        pixel_data[37][30] = 4'b1010; // x=30, y=37
        pixel_data[37][31] = 4'b0100; // x=31, y=37
        pixel_data[37][32] = 4'b1110; // x=32, y=37
        pixel_data[37][33] = 4'b0001; // x=33, y=37
        pixel_data[37][34] = 4'b1011; // x=34, y=37
        pixel_data[37][35] = 4'b0001; // x=35, y=37
        pixel_data[37][36] = 4'b0001; // x=36, y=37
        pixel_data[37][37] = 4'b0001; // x=37, y=37
        pixel_data[37][38] = 4'b0001; // x=38, y=37
        pixel_data[37][39] = 4'b0001; // x=39, y=37
        pixel_data[37][40] = 4'b0001; // x=40, y=37
        pixel_data[37][41] = 4'b0001; // x=41, y=37
        pixel_data[37][42] = 4'b0001; // x=42, y=37
        pixel_data[37][43] = 4'b0001; // x=43, y=37
        pixel_data[37][44] = 4'b0001; // x=44, y=37
        pixel_data[37][45] = 4'b0001; // x=45, y=37
        pixel_data[37][46] = 4'b0001; // x=46, y=37
        pixel_data[37][47] = 4'b0001; // x=47, y=37
        pixel_data[37][48] = 4'b0001; // x=48, y=37
        pixel_data[37][49] = 4'b0001; // x=49, y=37
        pixel_data[37][50] = 4'b0001; // x=50, y=37
        pixel_data[37][51] = 4'b0001; // x=51, y=37
        pixel_data[37][52] = 4'b0001; // x=52, y=37
        pixel_data[37][53] = 4'b0001; // x=53, y=37
        pixel_data[37][54] = 4'b0001; // x=54, y=37
        pixel_data[37][55] = 4'b0001; // x=55, y=37
        pixel_data[37][56] = 4'b0001; // x=56, y=37
        pixel_data[37][57] = 4'b0001; // x=57, y=37
        pixel_data[37][58] = 4'b0001; // x=58, y=37
        pixel_data[37][59] = 4'b0001; // x=59, y=37
        pixel_data[38][0] = 4'b0001; // x=0, y=38
        pixel_data[38][1] = 4'b0001; // x=1, y=38
        pixel_data[38][2] = 4'b0001; // x=2, y=38
        pixel_data[38][3] = 4'b0001; // x=3, y=38
        pixel_data[38][4] = 4'b0001; // x=4, y=38
        pixel_data[38][5] = 4'b0001; // x=5, y=38
        pixel_data[38][6] = 4'b0001; // x=6, y=38
        pixel_data[38][7] = 4'b0001; // x=7, y=38
        pixel_data[38][8] = 4'b0001; // x=8, y=38
        pixel_data[38][9] = 4'b0001; // x=9, y=38
        pixel_data[38][10] = 4'b0001; // x=10, y=38
        pixel_data[38][11] = 4'b0001; // x=11, y=38
        pixel_data[38][12] = 4'b0001; // x=12, y=38
        pixel_data[38][13] = 4'b0001; // x=13, y=38
        pixel_data[38][14] = 4'b0001; // x=14, y=38
        pixel_data[38][15] = 4'b0001; // x=15, y=38
        pixel_data[38][16] = 4'b0001; // x=16, y=38
        pixel_data[38][17] = 4'b0001; // x=17, y=38
        pixel_data[38][18] = 4'b0001; // x=18, y=38
        pixel_data[38][19] = 4'b0001; // x=19, y=38
        pixel_data[38][20] = 4'b0001; // x=20, y=38
        pixel_data[38][21] = 4'b0001; // x=21, y=38
        pixel_data[38][22] = 4'b0001; // x=22, y=38
        pixel_data[38][23] = 4'b0001; // x=23, y=38
        pixel_data[38][24] = 4'b0111; // x=24, y=38
        pixel_data[38][25] = 4'b1010; // x=25, y=38
        pixel_data[38][26] = 4'b0010; // x=26, y=38
        pixel_data[38][27] = 4'b0010; // x=27, y=38
        pixel_data[38][28] = 4'b1010; // x=28, y=38
        pixel_data[38][29] = 4'b0010; // x=29, y=38
        pixel_data[38][30] = 4'b1010; // x=30, y=38
        pixel_data[38][31] = 4'b1001; // x=31, y=38
        pixel_data[38][32] = 4'b0001; // x=32, y=38
        pixel_data[38][33] = 4'b1011; // x=33, y=38
        pixel_data[38][34] = 4'b0001; // x=34, y=38
        pixel_data[38][35] = 4'b0001; // x=35, y=38
        pixel_data[38][36] = 4'b0001; // x=36, y=38
        pixel_data[38][37] = 4'b0001; // x=37, y=38
        pixel_data[38][38] = 4'b0001; // x=38, y=38
        pixel_data[38][39] = 4'b0001; // x=39, y=38
        pixel_data[38][40] = 4'b0001; // x=40, y=38
        pixel_data[38][41] = 4'b0001; // x=41, y=38
        pixel_data[38][42] = 4'b0001; // x=42, y=38
        pixel_data[38][43] = 4'b0001; // x=43, y=38
        pixel_data[38][44] = 4'b0001; // x=44, y=38
        pixel_data[38][45] = 4'b0001; // x=45, y=38
        pixel_data[38][46] = 4'b0001; // x=46, y=38
        pixel_data[38][47] = 4'b0001; // x=47, y=38
        pixel_data[38][48] = 4'b0001; // x=48, y=38
        pixel_data[38][49] = 4'b0001; // x=49, y=38
        pixel_data[38][50] = 4'b0001; // x=50, y=38
        pixel_data[38][51] = 4'b0001; // x=51, y=38
        pixel_data[38][52] = 4'b0001; // x=52, y=38
        pixel_data[38][53] = 4'b0001; // x=53, y=38
        pixel_data[38][54] = 4'b0001; // x=54, y=38
        pixel_data[38][55] = 4'b0001; // x=55, y=38
        pixel_data[38][56] = 4'b0001; // x=56, y=38
        pixel_data[38][57] = 4'b0001; // x=57, y=38
        pixel_data[38][58] = 4'b0001; // x=58, y=38
        pixel_data[38][59] = 4'b0001; // x=59, y=38
        pixel_data[39][0] = 4'b0001; // x=0, y=39
        pixel_data[39][1] = 4'b0001; // x=1, y=39
        pixel_data[39][2] = 4'b0001; // x=2, y=39
        pixel_data[39][3] = 4'b0001; // x=3, y=39
        pixel_data[39][4] = 4'b0001; // x=4, y=39
        pixel_data[39][5] = 4'b0001; // x=5, y=39
        pixel_data[39][6] = 4'b0001; // x=6, y=39
        pixel_data[39][7] = 4'b0001; // x=7, y=39
        pixel_data[39][8] = 4'b0001; // x=8, y=39
        pixel_data[39][9] = 4'b0001; // x=9, y=39
        pixel_data[39][10] = 4'b0001; // x=10, y=39
        pixel_data[39][11] = 4'b0001; // x=11, y=39
        pixel_data[39][12] = 4'b0001; // x=12, y=39
        pixel_data[39][13] = 4'b0001; // x=13, y=39
        pixel_data[39][14] = 4'b0001; // x=14, y=39
        pixel_data[39][15] = 4'b0001; // x=15, y=39
        pixel_data[39][16] = 4'b0001; // x=16, y=39
        pixel_data[39][17] = 4'b0001; // x=17, y=39
        pixel_data[39][18] = 4'b0001; // x=18, y=39
        pixel_data[39][19] = 4'b1011; // x=19, y=39
        pixel_data[39][20] = 4'b0001; // x=20, y=39
        pixel_data[39][21] = 4'b1011; // x=21, y=39
        pixel_data[39][22] = 4'b0001; // x=22, y=39
        pixel_data[39][23] = 4'b1001; // x=23, y=39
        pixel_data[39][24] = 4'b1010; // x=24, y=39
        pixel_data[39][25] = 4'b0010; // x=25, y=39
        pixel_data[39][26] = 4'b0010; // x=26, y=39
        pixel_data[39][27] = 4'b1010; // x=27, y=39
        pixel_data[39][28] = 4'b0010; // x=28, y=39
        pixel_data[39][29] = 4'b1010; // x=29, y=39
        pixel_data[39][30] = 4'b0000; // x=30, y=39
        pixel_data[39][31] = 4'b1011; // x=31, y=39
        pixel_data[39][32] = 4'b1011; // x=32, y=39
        pixel_data[39][33] = 4'b0001; // x=33, y=39
        pixel_data[39][34] = 4'b0001; // x=34, y=39
        pixel_data[39][35] = 4'b0001; // x=35, y=39
        pixel_data[39][36] = 4'b0001; // x=36, y=39
        pixel_data[39][37] = 4'b0001; // x=37, y=39
        pixel_data[39][38] = 4'b0001; // x=38, y=39
        pixel_data[39][39] = 4'b0001; // x=39, y=39
        pixel_data[39][40] = 4'b0001; // x=40, y=39
        pixel_data[39][41] = 4'b0001; // x=41, y=39
        pixel_data[39][42] = 4'b0001; // x=42, y=39
        pixel_data[39][43] = 4'b0001; // x=43, y=39
        pixel_data[39][44] = 4'b0001; // x=44, y=39
        pixel_data[39][45] = 4'b0001; // x=45, y=39
        pixel_data[39][46] = 4'b0001; // x=46, y=39
        pixel_data[39][47] = 4'b0001; // x=47, y=39
        pixel_data[39][48] = 4'b0001; // x=48, y=39
        pixel_data[39][49] = 4'b0001; // x=49, y=39
        pixel_data[39][50] = 4'b0001; // x=50, y=39
        pixel_data[39][51] = 4'b0001; // x=51, y=39
        pixel_data[39][52] = 4'b0001; // x=52, y=39
        pixel_data[39][53] = 4'b0001; // x=53, y=39
        pixel_data[39][54] = 4'b0001; // x=54, y=39
        pixel_data[39][55] = 4'b0001; // x=55, y=39
        pixel_data[39][56] = 4'b0001; // x=56, y=39
        pixel_data[39][57] = 4'b0001; // x=57, y=39
        pixel_data[39][58] = 4'b0001; // x=58, y=39
        pixel_data[39][59] = 4'b0001; // x=59, y=39
        pixel_data[40][0] = 4'b0001; // x=0, y=40
        pixel_data[40][1] = 4'b0001; // x=1, y=40
        pixel_data[40][2] = 4'b0001; // x=2, y=40
        pixel_data[40][3] = 4'b0001; // x=3, y=40
        pixel_data[40][4] = 4'b0001; // x=4, y=40
        pixel_data[40][5] = 4'b0001; // x=5, y=40
        pixel_data[40][6] = 4'b0001; // x=6, y=40
        pixel_data[40][7] = 4'b0001; // x=7, y=40
        pixel_data[40][8] = 4'b0001; // x=8, y=40
        pixel_data[40][9] = 4'b0001; // x=9, y=40
        pixel_data[40][10] = 4'b0001; // x=10, y=40
        pixel_data[40][11] = 4'b0001; // x=11, y=40
        pixel_data[40][12] = 4'b0001; // x=12, y=40
        pixel_data[40][13] = 4'b0001; // x=13, y=40
        pixel_data[40][14] = 4'b0001; // x=14, y=40
        pixel_data[40][15] = 4'b0001; // x=15, y=40
        pixel_data[40][16] = 4'b0001; // x=16, y=40
        pixel_data[40][17] = 4'b0001; // x=17, y=40
        pixel_data[40][18] = 4'b0001; // x=18, y=40
        pixel_data[40][19] = 4'b1011; // x=19, y=40
        pixel_data[40][20] = 4'b1011; // x=20, y=40
        pixel_data[40][21] = 4'b0001; // x=21, y=40
        pixel_data[40][22] = 4'b1110; // x=22, y=40
        pixel_data[40][23] = 4'b0100; // x=23, y=40
        pixel_data[40][24] = 4'b1010; // x=24, y=40
        pixel_data[40][25] = 4'b0010; // x=25, y=40
        pixel_data[40][26] = 4'b0010; // x=26, y=40
        pixel_data[40][27] = 4'b0010; // x=27, y=40
        pixel_data[40][28] = 4'b0010; // x=28, y=40
        pixel_data[40][29] = 4'b1010; // x=29, y=40
        pixel_data[40][30] = 4'b1111; // x=30, y=40
        pixel_data[40][31] = 4'b0001; // x=31, y=40
        pixel_data[40][32] = 4'b1011; // x=32, y=40
        pixel_data[40][33] = 4'b0001; // x=33, y=40
        pixel_data[40][34] = 4'b0001; // x=34, y=40
        pixel_data[40][35] = 4'b0001; // x=35, y=40
        pixel_data[40][36] = 4'b0001; // x=36, y=40
        pixel_data[40][37] = 4'b0001; // x=37, y=40
        pixel_data[40][38] = 4'b0001; // x=38, y=40
        pixel_data[40][39] = 4'b0001; // x=39, y=40
        pixel_data[40][40] = 4'b0001; // x=40, y=40
        pixel_data[40][41] = 4'b0001; // x=41, y=40
        pixel_data[40][42] = 4'b0001; // x=42, y=40
        pixel_data[40][43] = 4'b0001; // x=43, y=40
        pixel_data[40][44] = 4'b0001; // x=44, y=40
        pixel_data[40][45] = 4'b0001; // x=45, y=40
        pixel_data[40][46] = 4'b0001; // x=46, y=40
        pixel_data[40][47] = 4'b0001; // x=47, y=40
        pixel_data[40][48] = 4'b0001; // x=48, y=40
        pixel_data[40][49] = 4'b0001; // x=49, y=40
        pixel_data[40][50] = 4'b0001; // x=50, y=40
        pixel_data[40][51] = 4'b0001; // x=51, y=40
        pixel_data[40][52] = 4'b0001; // x=52, y=40
        pixel_data[40][53] = 4'b0001; // x=53, y=40
        pixel_data[40][54] = 4'b0001; // x=54, y=40
        pixel_data[40][55] = 4'b0001; // x=55, y=40
        pixel_data[40][56] = 4'b0001; // x=56, y=40
        pixel_data[40][57] = 4'b0001; // x=57, y=40
        pixel_data[40][58] = 4'b0001; // x=58, y=40
        pixel_data[40][59] = 4'b0001; // x=59, y=40
        pixel_data[41][0] = 4'b0001; // x=0, y=41
        pixel_data[41][1] = 4'b0001; // x=1, y=41
        pixel_data[41][2] = 4'b0001; // x=2, y=41
        pixel_data[41][3] = 4'b0001; // x=3, y=41
        pixel_data[41][4] = 4'b0001; // x=4, y=41
        pixel_data[41][5] = 4'b0001; // x=5, y=41
        pixel_data[41][6] = 4'b0001; // x=6, y=41
        pixel_data[41][7] = 4'b0001; // x=7, y=41
        pixel_data[41][8] = 4'b0001; // x=8, y=41
        pixel_data[41][9] = 4'b0001; // x=9, y=41
        pixel_data[41][10] = 4'b0001; // x=10, y=41
        pixel_data[41][11] = 4'b0001; // x=11, y=41
        pixel_data[41][12] = 4'b0001; // x=12, y=41
        pixel_data[41][13] = 4'b0001; // x=13, y=41
        pixel_data[41][14] = 4'b0001; // x=14, y=41
        pixel_data[41][15] = 4'b0001; // x=15, y=41
        pixel_data[41][16] = 4'b0001; // x=16, y=41
        pixel_data[41][17] = 4'b0001; // x=17, y=41
        pixel_data[41][18] = 4'b0001; // x=18, y=41
        pixel_data[41][19] = 4'b0001; // x=19, y=41
        pixel_data[41][20] = 4'b1011; // x=20, y=41
        pixel_data[41][21] = 4'b0001; // x=21, y=41
        pixel_data[41][22] = 4'b0101; // x=22, y=41
        pixel_data[41][23] = 4'b1010; // x=23, y=41
        pixel_data[41][24] = 4'b0010; // x=24, y=41
        pixel_data[41][25] = 4'b1010; // x=25, y=41
        pixel_data[41][26] = 4'b1010; // x=26, y=41
        pixel_data[41][27] = 4'b0010; // x=27, y=41
        pixel_data[41][28] = 4'b1010; // x=28, y=41
        pixel_data[41][29] = 4'b1101; // x=29, y=41
        pixel_data[41][30] = 4'b0001; // x=30, y=41
        pixel_data[41][31] = 4'b1011; // x=31, y=41
        pixel_data[41][32] = 4'b0001; // x=32, y=41
        pixel_data[41][33] = 4'b0001; // x=33, y=41
        pixel_data[41][34] = 4'b0001; // x=34, y=41
        pixel_data[41][35] = 4'b0001; // x=35, y=41
        pixel_data[41][36] = 4'b0001; // x=36, y=41
        pixel_data[41][37] = 4'b0001; // x=37, y=41
        pixel_data[41][38] = 4'b0001; // x=38, y=41
        pixel_data[41][39] = 4'b0001; // x=39, y=41
        pixel_data[41][40] = 4'b0001; // x=40, y=41
        pixel_data[41][41] = 4'b0001; // x=41, y=41
        pixel_data[41][42] = 4'b0001; // x=42, y=41
        pixel_data[41][43] = 4'b0001; // x=43, y=41
        pixel_data[41][44] = 4'b0001; // x=44, y=41
        pixel_data[41][45] = 4'b0001; // x=45, y=41
        pixel_data[41][46] = 4'b0001; // x=46, y=41
        pixel_data[41][47] = 4'b0001; // x=47, y=41
        pixel_data[41][48] = 4'b0001; // x=48, y=41
        pixel_data[41][49] = 4'b0001; // x=49, y=41
        pixel_data[41][50] = 4'b0001; // x=50, y=41
        pixel_data[41][51] = 4'b0001; // x=51, y=41
        pixel_data[41][52] = 4'b0001; // x=52, y=41
        pixel_data[41][53] = 4'b0001; // x=53, y=41
        pixel_data[41][54] = 4'b0001; // x=54, y=41
        pixel_data[41][55] = 4'b0001; // x=55, y=41
        pixel_data[41][56] = 4'b0001; // x=56, y=41
        pixel_data[41][57] = 4'b0001; // x=57, y=41
        pixel_data[41][58] = 4'b0001; // x=58, y=41
        pixel_data[41][59] = 4'b0001; // x=59, y=41
        pixel_data[42][0] = 4'b0001; // x=0, y=42
        pixel_data[42][1] = 4'b0001; // x=1, y=42
        pixel_data[42][2] = 4'b0001; // x=2, y=42
        pixel_data[42][3] = 4'b0001; // x=3, y=42
        pixel_data[42][4] = 4'b0001; // x=4, y=42
        pixel_data[42][5] = 4'b0001; // x=5, y=42
        pixel_data[42][6] = 4'b0001; // x=6, y=42
        pixel_data[42][7] = 4'b0001; // x=7, y=42
        pixel_data[42][8] = 4'b0001; // x=8, y=42
        pixel_data[42][9] = 4'b0001; // x=9, y=42
        pixel_data[42][10] = 4'b0001; // x=10, y=42
        pixel_data[42][11] = 4'b0001; // x=11, y=42
        pixel_data[42][12] = 4'b0001; // x=12, y=42
        pixel_data[42][13] = 4'b0001; // x=13, y=42
        pixel_data[42][14] = 4'b0001; // x=14, y=42
        pixel_data[42][15] = 4'b0001; // x=15, y=42
        pixel_data[42][16] = 4'b0001; // x=16, y=42
        pixel_data[42][17] = 4'b0001; // x=17, y=42
        pixel_data[42][18] = 4'b0001; // x=18, y=42
        pixel_data[42][19] = 4'b1011; // x=19, y=42
        pixel_data[42][20] = 4'b0001; // x=20, y=42
        pixel_data[42][21] = 4'b0110; // x=21, y=42
        pixel_data[42][22] = 4'b0010; // x=22, y=42
        pixel_data[42][23] = 4'b0010; // x=23, y=42
        pixel_data[42][24] = 4'b0010; // x=24, y=42
        pixel_data[42][25] = 4'b0010; // x=25, y=42
        pixel_data[42][26] = 4'b0010; // x=26, y=42
        pixel_data[42][27] = 4'b0010; // x=27, y=42
        pixel_data[42][28] = 4'b0100; // x=28, y=42
        pixel_data[42][29] = 4'b0110; // x=29, y=42
        pixel_data[42][30] = 4'b0001; // x=30, y=42
        pixel_data[42][31] = 4'b1011; // x=31, y=42
        pixel_data[42][32] = 4'b0001; // x=32, y=42
        pixel_data[42][33] = 4'b0001; // x=33, y=42
        pixel_data[42][34] = 4'b0001; // x=34, y=42
        pixel_data[42][35] = 4'b0001; // x=35, y=42
        pixel_data[42][36] = 4'b0001; // x=36, y=42
        pixel_data[42][37] = 4'b0001; // x=37, y=42
        pixel_data[42][38] = 4'b0001; // x=38, y=42
        pixel_data[42][39] = 4'b0001; // x=39, y=42
        pixel_data[42][40] = 4'b0001; // x=40, y=42
        pixel_data[42][41] = 4'b0001; // x=41, y=42
        pixel_data[42][42] = 4'b0001; // x=42, y=42
        pixel_data[42][43] = 4'b0001; // x=43, y=42
        pixel_data[42][44] = 4'b0001; // x=44, y=42
        pixel_data[42][45] = 4'b0001; // x=45, y=42
        pixel_data[42][46] = 4'b0001; // x=46, y=42
        pixel_data[42][47] = 4'b0001; // x=47, y=42
        pixel_data[42][48] = 4'b0001; // x=48, y=42
        pixel_data[42][49] = 4'b0001; // x=49, y=42
        pixel_data[42][50] = 4'b0001; // x=50, y=42
        pixel_data[42][51] = 4'b0001; // x=51, y=42
        pixel_data[42][52] = 4'b0001; // x=52, y=42
        pixel_data[42][53] = 4'b0001; // x=53, y=42
        pixel_data[42][54] = 4'b0001; // x=54, y=42
        pixel_data[42][55] = 4'b0001; // x=55, y=42
        pixel_data[42][56] = 4'b0001; // x=56, y=42
        pixel_data[42][57] = 4'b0001; // x=57, y=42
        pixel_data[42][58] = 4'b0001; // x=58, y=42
        pixel_data[42][59] = 4'b0001; // x=59, y=42
        pixel_data[43][0] = 4'b0001; // x=0, y=43
        pixel_data[43][1] = 4'b0001; // x=1, y=43
        pixel_data[43][2] = 4'b0001; // x=2, y=43
        pixel_data[43][3] = 4'b0001; // x=3, y=43
        pixel_data[43][4] = 4'b0001; // x=4, y=43
        pixel_data[43][5] = 4'b0001; // x=5, y=43
        pixel_data[43][6] = 4'b0001; // x=6, y=43
        pixel_data[43][7] = 4'b0001; // x=7, y=43
        pixel_data[43][8] = 4'b0001; // x=8, y=43
        pixel_data[43][9] = 4'b0001; // x=9, y=43
        pixel_data[43][10] = 4'b0001; // x=10, y=43
        pixel_data[43][11] = 4'b0001; // x=11, y=43
        pixel_data[43][12] = 4'b0001; // x=12, y=43
        pixel_data[43][13] = 4'b0001; // x=13, y=43
        pixel_data[43][14] = 4'b0001; // x=14, y=43
        pixel_data[43][15] = 4'b0001; // x=15, y=43
        pixel_data[43][16] = 4'b0001; // x=16, y=43
        pixel_data[43][17] = 4'b0001; // x=17, y=43
        pixel_data[43][18] = 4'b0001; // x=18, y=43
        pixel_data[43][19] = 4'b1011; // x=19, y=43
        pixel_data[43][20] = 4'b1011; // x=20, y=43
        pixel_data[43][21] = 4'b0111; // x=21, y=43
        pixel_data[43][22] = 4'b1010; // x=22, y=43
        pixel_data[43][23] = 4'b0010; // x=23, y=43
        pixel_data[43][24] = 4'b1010; // x=24, y=43
        pixel_data[43][25] = 4'b1010; // x=25, y=43
        pixel_data[43][26] = 4'b0010; // x=26, y=43
        pixel_data[43][27] = 4'b1010; // x=27, y=43
        pixel_data[43][28] = 4'b1100; // x=28, y=43
        pixel_data[43][29] = 4'b0001; // x=29, y=43
        pixel_data[43][30] = 4'b1011; // x=30, y=43
        pixel_data[43][31] = 4'b0001; // x=31, y=43
        pixel_data[43][32] = 4'b0001; // x=32, y=43
        pixel_data[43][33] = 4'b0001; // x=33, y=43
        pixel_data[43][34] = 4'b0001; // x=34, y=43
        pixel_data[43][35] = 4'b0001; // x=35, y=43
        pixel_data[43][36] = 4'b0001; // x=36, y=43
        pixel_data[43][37] = 4'b0001; // x=37, y=43
        pixel_data[43][38] = 4'b0001; // x=38, y=43
        pixel_data[43][39] = 4'b0001; // x=39, y=43
        pixel_data[43][40] = 4'b0001; // x=40, y=43
        pixel_data[43][41] = 4'b0001; // x=41, y=43
        pixel_data[43][42] = 4'b0001; // x=42, y=43
        pixel_data[43][43] = 4'b0001; // x=43, y=43
        pixel_data[43][44] = 4'b0001; // x=44, y=43
        pixel_data[43][45] = 4'b0001; // x=45, y=43
        pixel_data[43][46] = 4'b0001; // x=46, y=43
        pixel_data[43][47] = 4'b0001; // x=47, y=43
        pixel_data[43][48] = 4'b0001; // x=48, y=43
        pixel_data[43][49] = 4'b0001; // x=49, y=43
        pixel_data[43][50] = 4'b0001; // x=50, y=43
        pixel_data[43][51] = 4'b0001; // x=51, y=43
        pixel_data[43][52] = 4'b0001; // x=52, y=43
        pixel_data[43][53] = 4'b0001; // x=53, y=43
        pixel_data[43][54] = 4'b0001; // x=54, y=43
        pixel_data[43][55] = 4'b0001; // x=55, y=43
        pixel_data[43][56] = 4'b0001; // x=56, y=43
        pixel_data[43][57] = 4'b0001; // x=57, y=43
        pixel_data[43][58] = 4'b0001; // x=58, y=43
        pixel_data[43][59] = 4'b0001; // x=59, y=43
        pixel_data[44][0] = 4'b0001; // x=0, y=44
        pixel_data[44][1] = 4'b0001; // x=1, y=44
        pixel_data[44][2] = 4'b0001; // x=2, y=44
        pixel_data[44][3] = 4'b0001; // x=3, y=44
        pixel_data[44][4] = 4'b0001; // x=4, y=44
        pixel_data[44][5] = 4'b0001; // x=5, y=44
        pixel_data[44][6] = 4'b0001; // x=6, y=44
        pixel_data[44][7] = 4'b0001; // x=7, y=44
        pixel_data[44][8] = 4'b0001; // x=8, y=44
        pixel_data[44][9] = 4'b0001; // x=9, y=44
        pixel_data[44][10] = 4'b0001; // x=10, y=44
        pixel_data[44][11] = 4'b0001; // x=11, y=44
        pixel_data[44][12] = 4'b0001; // x=12, y=44
        pixel_data[44][13] = 4'b0001; // x=13, y=44
        pixel_data[44][14] = 4'b0001; // x=14, y=44
        pixel_data[44][15] = 4'b0001; // x=15, y=44
        pixel_data[44][16] = 4'b0001; // x=16, y=44
        pixel_data[44][17] = 4'b0001; // x=17, y=44
        pixel_data[44][18] = 4'b0001; // x=18, y=44
        pixel_data[44][19] = 4'b0001; // x=19, y=44
        pixel_data[44][20] = 4'b1001; // x=20, y=44
        pixel_data[44][21] = 4'b1010; // x=21, y=44
        pixel_data[44][22] = 4'b0010; // x=22, y=44
        pixel_data[44][23] = 4'b0010; // x=23, y=44
        pixel_data[44][24] = 4'b0010; // x=24, y=44
        pixel_data[44][25] = 4'b0010; // x=25, y=44
        pixel_data[44][26] = 4'b0010; // x=26, y=44
        pixel_data[44][27] = 4'b0100; // x=27, y=44
        pixel_data[44][28] = 4'b1000; // x=28, y=44
        pixel_data[44][29] = 4'b0001; // x=29, y=44
        pixel_data[44][30] = 4'b1011; // x=30, y=44
        pixel_data[44][31] = 4'b0001; // x=31, y=44
        pixel_data[44][32] = 4'b0001; // x=32, y=44
        pixel_data[44][33] = 4'b0001; // x=33, y=44
        pixel_data[44][34] = 4'b0001; // x=34, y=44
        pixel_data[44][35] = 4'b0001; // x=35, y=44
        pixel_data[44][36] = 4'b0001; // x=36, y=44
        pixel_data[44][37] = 4'b0001; // x=37, y=44
        pixel_data[44][38] = 4'b0001; // x=38, y=44
        pixel_data[44][39] = 4'b0001; // x=39, y=44
        pixel_data[44][40] = 4'b0001; // x=40, y=44
        pixel_data[44][41] = 4'b0001; // x=41, y=44
        pixel_data[44][42] = 4'b0001; // x=42, y=44
        pixel_data[44][43] = 4'b0001; // x=43, y=44
        pixel_data[44][44] = 4'b0001; // x=44, y=44
        pixel_data[44][45] = 4'b0001; // x=45, y=44
        pixel_data[44][46] = 4'b0001; // x=46, y=44
        pixel_data[44][47] = 4'b0001; // x=47, y=44
        pixel_data[44][48] = 4'b0001; // x=48, y=44
        pixel_data[44][49] = 4'b0001; // x=49, y=44
        pixel_data[44][50] = 4'b0001; // x=50, y=44
        pixel_data[44][51] = 4'b0001; // x=51, y=44
        pixel_data[44][52] = 4'b0001; // x=52, y=44
        pixel_data[44][53] = 4'b0001; // x=53, y=44
        pixel_data[44][54] = 4'b0001; // x=54, y=44
        pixel_data[44][55] = 4'b0001; // x=55, y=44
        pixel_data[44][56] = 4'b0001; // x=56, y=44
        pixel_data[44][57] = 4'b0001; // x=57, y=44
        pixel_data[44][58] = 4'b0001; // x=58, y=44
        pixel_data[44][59] = 4'b0001; // x=59, y=44
        pixel_data[45][0] = 4'b0001; // x=0, y=45
        pixel_data[45][1] = 4'b0001; // x=1, y=45
        pixel_data[45][2] = 4'b0001; // x=2, y=45
        pixel_data[45][3] = 4'b0001; // x=3, y=45
        pixel_data[45][4] = 4'b0001; // x=4, y=45
        pixel_data[45][5] = 4'b0001; // x=5, y=45
        pixel_data[45][6] = 4'b0001; // x=6, y=45
        pixel_data[45][7] = 4'b0001; // x=7, y=45
        pixel_data[45][8] = 4'b0001; // x=8, y=45
        pixel_data[45][9] = 4'b0001; // x=9, y=45
        pixel_data[45][10] = 4'b0001; // x=10, y=45
        pixel_data[45][11] = 4'b0001; // x=11, y=45
        pixel_data[45][12] = 4'b0001; // x=12, y=45
        pixel_data[45][13] = 4'b0001; // x=13, y=45
        pixel_data[45][14] = 4'b0001; // x=14, y=45
        pixel_data[45][15] = 4'b0001; // x=15, y=45
        pixel_data[45][16] = 4'b0001; // x=16, y=45
        pixel_data[45][17] = 4'b0001; // x=17, y=45
        pixel_data[45][18] = 4'b0001; // x=18, y=45
        pixel_data[45][19] = 4'b1110; // x=19, y=45
        pixel_data[45][20] = 4'b0010; // x=20, y=45
        pixel_data[45][21] = 4'b1010; // x=21, y=45
        pixel_data[45][22] = 4'b1010; // x=22, y=45
        pixel_data[45][23] = 4'b1010; // x=23, y=45
        pixel_data[45][24] = 4'b1010; // x=24, y=45
        pixel_data[45][25] = 4'b1010; // x=25, y=45
        pixel_data[45][26] = 4'b1010; // x=26, y=45
        pixel_data[45][27] = 4'b0011; // x=27, y=45
        pixel_data[45][28] = 4'b0001; // x=28, y=45
        pixel_data[45][29] = 4'b1011; // x=29, y=45
        pixel_data[45][30] = 4'b1011; // x=30, y=45
        pixel_data[45][31] = 4'b1011; // x=31, y=45
        pixel_data[45][32] = 4'b0001; // x=32, y=45
        pixel_data[45][33] = 4'b0001; // x=33, y=45
        pixel_data[45][34] = 4'b0001; // x=34, y=45
        pixel_data[45][35] = 4'b0001; // x=35, y=45
        pixel_data[45][36] = 4'b0001; // x=36, y=45
        pixel_data[45][37] = 4'b0001; // x=37, y=45
        pixel_data[45][38] = 4'b0001; // x=38, y=45
        pixel_data[45][39] = 4'b0001; // x=39, y=45
        pixel_data[45][40] = 4'b0001; // x=40, y=45
        pixel_data[45][41] = 4'b0001; // x=41, y=45
        pixel_data[45][42] = 4'b0001; // x=42, y=45
        pixel_data[45][43] = 4'b0001; // x=43, y=45
        pixel_data[45][44] = 4'b0001; // x=44, y=45
        pixel_data[45][45] = 4'b0001; // x=45, y=45
        pixel_data[45][46] = 4'b0001; // x=46, y=45
        pixel_data[45][47] = 4'b0001; // x=47, y=45
        pixel_data[45][48] = 4'b0001; // x=48, y=45
        pixel_data[45][49] = 4'b0001; // x=49, y=45
        pixel_data[45][50] = 4'b0001; // x=50, y=45
        pixel_data[45][51] = 4'b0001; // x=51, y=45
        pixel_data[45][52] = 4'b0001; // x=52, y=45
        pixel_data[45][53] = 4'b0001; // x=53, y=45
        pixel_data[45][54] = 4'b0001; // x=54, y=45
        pixel_data[45][55] = 4'b0001; // x=55, y=45
        pixel_data[45][56] = 4'b0001; // x=56, y=45
        pixel_data[45][57] = 4'b0001; // x=57, y=45
        pixel_data[45][58] = 4'b0001; // x=58, y=45
        pixel_data[45][59] = 4'b0001; // x=59, y=45
        pixel_data[46][0] = 4'b0001; // x=0, y=46
        pixel_data[46][1] = 4'b0001; // x=1, y=46
        pixel_data[46][2] = 4'b0001; // x=2, y=46
        pixel_data[46][3] = 4'b0001; // x=3, y=46
        pixel_data[46][4] = 4'b0001; // x=4, y=46
        pixel_data[46][5] = 4'b0001; // x=5, y=46
        pixel_data[46][6] = 4'b0001; // x=6, y=46
        pixel_data[46][7] = 4'b0001; // x=7, y=46
        pixel_data[46][8] = 4'b0001; // x=8, y=46
        pixel_data[46][9] = 4'b0001; // x=9, y=46
        pixel_data[46][10] = 4'b0001; // x=10, y=46
        pixel_data[46][11] = 4'b0001; // x=11, y=46
        pixel_data[46][12] = 4'b0001; // x=12, y=46
        pixel_data[46][13] = 4'b0001; // x=13, y=46
        pixel_data[46][14] = 4'b0001; // x=14, y=46
        pixel_data[46][15] = 4'b0001; // x=15, y=46
        pixel_data[46][16] = 4'b0001; // x=16, y=46
        pixel_data[46][17] = 4'b1011; // x=17, y=46
        pixel_data[46][18] = 4'b0001; // x=18, y=46
        pixel_data[46][19] = 4'b1001; // x=19, y=46
        pixel_data[46][20] = 4'b0000; // x=20, y=46
        pixel_data[46][21] = 4'b0111; // x=21, y=46
        pixel_data[46][22] = 4'b0111; // x=22, y=46
        pixel_data[46][23] = 4'b0111; // x=23, y=46
        pixel_data[46][24] = 4'b0111; // x=24, y=46
        pixel_data[46][25] = 4'b0000; // x=25, y=46
        pixel_data[46][26] = 4'b0101; // x=26, y=46
        pixel_data[46][27] = 4'b1011; // x=27, y=46
        pixel_data[46][28] = 4'b0001; // x=28, y=46
        pixel_data[46][29] = 4'b0001; // x=29, y=46
        pixel_data[46][30] = 4'b0001; // x=30, y=46
        pixel_data[46][31] = 4'b0001; // x=31, y=46
        pixel_data[46][32] = 4'b0001; // x=32, y=46
        pixel_data[46][33] = 4'b0001; // x=33, y=46
        pixel_data[46][34] = 4'b0001; // x=34, y=46
        pixel_data[46][35] = 4'b0001; // x=35, y=46
        pixel_data[46][36] = 4'b0001; // x=36, y=46
        pixel_data[46][37] = 4'b0001; // x=37, y=46
        pixel_data[46][38] = 4'b0001; // x=38, y=46
        pixel_data[46][39] = 4'b0001; // x=39, y=46
        pixel_data[46][40] = 4'b0001; // x=40, y=46
        pixel_data[46][41] = 4'b0001; // x=41, y=46
        pixel_data[46][42] = 4'b0001; // x=42, y=46
        pixel_data[46][43] = 4'b0001; // x=43, y=46
        pixel_data[46][44] = 4'b0001; // x=44, y=46
        pixel_data[46][45] = 4'b0001; // x=45, y=46
        pixel_data[46][46] = 4'b0001; // x=46, y=46
        pixel_data[46][47] = 4'b0001; // x=47, y=46
        pixel_data[46][48] = 4'b0001; // x=48, y=46
        pixel_data[46][49] = 4'b0001; // x=49, y=46
        pixel_data[46][50] = 4'b0001; // x=50, y=46
        pixel_data[46][51] = 4'b0001; // x=51, y=46
        pixel_data[46][52] = 4'b0001; // x=52, y=46
        pixel_data[46][53] = 4'b0001; // x=53, y=46
        pixel_data[46][54] = 4'b0001; // x=54, y=46
        pixel_data[46][55] = 4'b0001; // x=55, y=46
        pixel_data[46][56] = 4'b0001; // x=56, y=46
        pixel_data[46][57] = 4'b0001; // x=57, y=46
        pixel_data[46][58] = 4'b0001; // x=58, y=46
        pixel_data[46][59] = 4'b0001; // x=59, y=46
        pixel_data[47][0] = 4'b0001; // x=0, y=47
        pixel_data[47][1] = 4'b0001; // x=1, y=47
        pixel_data[47][2] = 4'b0001; // x=2, y=47
        pixel_data[47][3] = 4'b0001; // x=3, y=47
        pixel_data[47][4] = 4'b0001; // x=4, y=47
        pixel_data[47][5] = 4'b0001; // x=5, y=47
        pixel_data[47][6] = 4'b0001; // x=6, y=47
        pixel_data[47][7] = 4'b0001; // x=7, y=47
        pixel_data[47][8] = 4'b0001; // x=8, y=47
        pixel_data[47][9] = 4'b0001; // x=9, y=47
        pixel_data[47][10] = 4'b0001; // x=10, y=47
        pixel_data[47][11] = 4'b0001; // x=11, y=47
        pixel_data[47][12] = 4'b0001; // x=12, y=47
        pixel_data[47][13] = 4'b0001; // x=13, y=47
        pixel_data[47][14] = 4'b0001; // x=14, y=47
        pixel_data[47][15] = 4'b0001; // x=15, y=47
        pixel_data[47][16] = 4'b0001; // x=16, y=47
        pixel_data[47][17] = 4'b0001; // x=17, y=47
        pixel_data[47][18] = 4'b0001; // x=18, y=47
        pixel_data[47][19] = 4'b0001; // x=19, y=47
        pixel_data[47][20] = 4'b0001; // x=20, y=47
        pixel_data[47][21] = 4'b0001; // x=21, y=47
        pixel_data[47][22] = 4'b0001; // x=22, y=47
        pixel_data[47][23] = 4'b0001; // x=23, y=47
        pixel_data[47][24] = 4'b0001; // x=24, y=47
        pixel_data[47][25] = 4'b0001; // x=25, y=47
        pixel_data[47][26] = 4'b0001; // x=26, y=47
        pixel_data[47][27] = 4'b1011; // x=27, y=47
        pixel_data[47][28] = 4'b0001; // x=28, y=47
        pixel_data[47][29] = 4'b0001; // x=29, y=47
        pixel_data[47][30] = 4'b0001; // x=30, y=47
        pixel_data[47][31] = 4'b0001; // x=31, y=47
        pixel_data[47][32] = 4'b0001; // x=32, y=47
        pixel_data[47][33] = 4'b0001; // x=33, y=47
        pixel_data[47][34] = 4'b0001; // x=34, y=47
        pixel_data[47][35] = 4'b0001; // x=35, y=47
        pixel_data[47][36] = 4'b0001; // x=36, y=47
        pixel_data[47][37] = 4'b0001; // x=37, y=47
        pixel_data[47][38] = 4'b0001; // x=38, y=47
        pixel_data[47][39] = 4'b0001; // x=39, y=47
        pixel_data[47][40] = 4'b0001; // x=40, y=47
        pixel_data[47][41] = 4'b0001; // x=41, y=47
        pixel_data[47][42] = 4'b0001; // x=42, y=47
        pixel_data[47][43] = 4'b0001; // x=43, y=47
        pixel_data[47][44] = 4'b0001; // x=44, y=47
        pixel_data[47][45] = 4'b0001; // x=45, y=47
        pixel_data[47][46] = 4'b0001; // x=46, y=47
        pixel_data[47][47] = 4'b0001; // x=47, y=47
        pixel_data[47][48] = 4'b0001; // x=48, y=47
        pixel_data[47][49] = 4'b0001; // x=49, y=47
        pixel_data[47][50] = 4'b0001; // x=50, y=47
        pixel_data[47][51] = 4'b0001; // x=51, y=47
        pixel_data[47][52] = 4'b0001; // x=52, y=47
        pixel_data[47][53] = 4'b0001; // x=53, y=47
        pixel_data[47][54] = 4'b0001; // x=54, y=47
        pixel_data[47][55] = 4'b0001; // x=55, y=47
        pixel_data[47][56] = 4'b0001; // x=56, y=47
        pixel_data[47][57] = 4'b0001; // x=57, y=47
        pixel_data[47][58] = 4'b0001; // x=58, y=47
        pixel_data[47][59] = 4'b0001; // x=59, y=47
        pixel_data[48][0] = 4'b0001; // x=0, y=48
        pixel_data[48][1] = 4'b0001; // x=1, y=48
        pixel_data[48][2] = 4'b0001; // x=2, y=48
        pixel_data[48][3] = 4'b0001; // x=3, y=48
        pixel_data[48][4] = 4'b0001; // x=4, y=48
        pixel_data[48][5] = 4'b0001; // x=5, y=48
        pixel_data[48][6] = 4'b0001; // x=6, y=48
        pixel_data[48][7] = 4'b0001; // x=7, y=48
        pixel_data[48][8] = 4'b0001; // x=8, y=48
        pixel_data[48][9] = 4'b0001; // x=9, y=48
        pixel_data[48][10] = 4'b0001; // x=10, y=48
        pixel_data[48][11] = 4'b0001; // x=11, y=48
        pixel_data[48][12] = 4'b0001; // x=12, y=48
        pixel_data[48][13] = 4'b0001; // x=13, y=48
        pixel_data[48][14] = 4'b0001; // x=14, y=48
        pixel_data[48][15] = 4'b0001; // x=15, y=48
        pixel_data[48][16] = 4'b0001; // x=16, y=48
        pixel_data[48][17] = 4'b0001; // x=17, y=48
        pixel_data[48][18] = 4'b1011; // x=18, y=48
        pixel_data[48][19] = 4'b1011; // x=19, y=48
        pixel_data[48][20] = 4'b1011; // x=20, y=48
        pixel_data[48][21] = 4'b1011; // x=21, y=48
        pixel_data[48][22] = 4'b1011; // x=22, y=48
        pixel_data[48][23] = 4'b1011; // x=23, y=48
        pixel_data[48][24] = 4'b1011; // x=24, y=48
        pixel_data[48][25] = 4'b1011; // x=25, y=48
        pixel_data[48][26] = 4'b1011; // x=26, y=48
        pixel_data[48][27] = 4'b0001; // x=27, y=48
        pixel_data[48][28] = 4'b0001; // x=28, y=48
        pixel_data[48][29] = 4'b0001; // x=29, y=48
        pixel_data[48][30] = 4'b0001; // x=30, y=48
        pixel_data[48][31] = 4'b0001; // x=31, y=48
        pixel_data[48][32] = 4'b0001; // x=32, y=48
        pixel_data[48][33] = 4'b0001; // x=33, y=48
        pixel_data[48][34] = 4'b0001; // x=34, y=48
        pixel_data[48][35] = 4'b0001; // x=35, y=48
        pixel_data[48][36] = 4'b0001; // x=36, y=48
        pixel_data[48][37] = 4'b0001; // x=37, y=48
        pixel_data[48][38] = 4'b0001; // x=38, y=48
        pixel_data[48][39] = 4'b0001; // x=39, y=48
        pixel_data[48][40] = 4'b0001; // x=40, y=48
        pixel_data[48][41] = 4'b0001; // x=41, y=48
        pixel_data[48][42] = 4'b0001; // x=42, y=48
        pixel_data[48][43] = 4'b0001; // x=43, y=48
        pixel_data[48][44] = 4'b0001; // x=44, y=48
        pixel_data[48][45] = 4'b0001; // x=45, y=48
        pixel_data[48][46] = 4'b0001; // x=46, y=48
        pixel_data[48][47] = 4'b0001; // x=47, y=48
        pixel_data[48][48] = 4'b0001; // x=48, y=48
        pixel_data[48][49] = 4'b0001; // x=49, y=48
        pixel_data[48][50] = 4'b0001; // x=50, y=48
        pixel_data[48][51] = 4'b0001; // x=51, y=48
        pixel_data[48][52] = 4'b0001; // x=52, y=48
        pixel_data[48][53] = 4'b0001; // x=53, y=48
        pixel_data[48][54] = 4'b0001; // x=54, y=48
        pixel_data[48][55] = 4'b0001; // x=55, y=48
        pixel_data[48][56] = 4'b0001; // x=56, y=48
        pixel_data[48][57] = 4'b0001; // x=57, y=48
        pixel_data[48][58] = 4'b0001; // x=58, y=48
        pixel_data[48][59] = 4'b0001; // x=59, y=48
        pixel_data[49][0] = 4'b0001; // x=0, y=49
        pixel_data[49][1] = 4'b0001; // x=1, y=49
        pixel_data[49][2] = 4'b0001; // x=2, y=49
        pixel_data[49][3] = 4'b0001; // x=3, y=49
        pixel_data[49][4] = 4'b0001; // x=4, y=49
        pixel_data[49][5] = 4'b0001; // x=5, y=49
        pixel_data[49][6] = 4'b0001; // x=6, y=49
        pixel_data[49][7] = 4'b0001; // x=7, y=49
        pixel_data[49][8] = 4'b0001; // x=8, y=49
        pixel_data[49][9] = 4'b0001; // x=9, y=49
        pixel_data[49][10] = 4'b0001; // x=10, y=49
        pixel_data[49][11] = 4'b0001; // x=11, y=49
        pixel_data[49][12] = 4'b0001; // x=12, y=49
        pixel_data[49][13] = 4'b0001; // x=13, y=49
        pixel_data[49][14] = 4'b0001; // x=14, y=49
        pixel_data[49][15] = 4'b0001; // x=15, y=49
        pixel_data[49][16] = 4'b0001; // x=16, y=49
        pixel_data[49][17] = 4'b0001; // x=17, y=49
        pixel_data[49][18] = 4'b0001; // x=18, y=49
        pixel_data[49][19] = 4'b0001; // x=19, y=49
        pixel_data[49][20] = 4'b0001; // x=20, y=49
        pixel_data[49][21] = 4'b0001; // x=21, y=49
        pixel_data[49][22] = 4'b0001; // x=22, y=49
        pixel_data[49][23] = 4'b0001; // x=23, y=49
        pixel_data[49][24] = 4'b0001; // x=24, y=49
        pixel_data[49][25] = 4'b0001; // x=25, y=49
        pixel_data[49][26] = 4'b0001; // x=26, y=49
        pixel_data[49][27] = 4'b0001; // x=27, y=49
        pixel_data[49][28] = 4'b0001; // x=28, y=49
        pixel_data[49][29] = 4'b0001; // x=29, y=49
        pixel_data[49][30] = 4'b0001; // x=30, y=49
        pixel_data[49][31] = 4'b0001; // x=31, y=49
        pixel_data[49][32] = 4'b0001; // x=32, y=49
        pixel_data[49][33] = 4'b0001; // x=33, y=49
        pixel_data[49][34] = 4'b0001; // x=34, y=49
        pixel_data[49][35] = 4'b0001; // x=35, y=49
        pixel_data[49][36] = 4'b0001; // x=36, y=49
        pixel_data[49][37] = 4'b0001; // x=37, y=49
        pixel_data[49][38] = 4'b0001; // x=38, y=49
        pixel_data[49][39] = 4'b0001; // x=39, y=49
        pixel_data[49][40] = 4'b0001; // x=40, y=49
        pixel_data[49][41] = 4'b0001; // x=41, y=49
        pixel_data[49][42] = 4'b0001; // x=42, y=49
        pixel_data[49][43] = 4'b0001; // x=43, y=49
        pixel_data[49][44] = 4'b0001; // x=44, y=49
        pixel_data[49][45] = 4'b0001; // x=45, y=49
        pixel_data[49][46] = 4'b0001; // x=46, y=49
        pixel_data[49][47] = 4'b0001; // x=47, y=49
        pixel_data[49][48] = 4'b0001; // x=48, y=49
        pixel_data[49][49] = 4'b0001; // x=49, y=49
        pixel_data[49][50] = 4'b0001; // x=50, y=49
        pixel_data[49][51] = 4'b0001; // x=51, y=49
        pixel_data[49][52] = 4'b0001; // x=52, y=49
        pixel_data[49][53] = 4'b0001; // x=53, y=49
        pixel_data[49][54] = 4'b0001; // x=54, y=49
        pixel_data[49][55] = 4'b0001; // x=55, y=49
        pixel_data[49][56] = 4'b0001; // x=56, y=49
        pixel_data[49][57] = 4'b0001; // x=57, y=49
        pixel_data[49][58] = 4'b0001; // x=58, y=49
        pixel_data[49][59] = 4'b0001; // x=59, y=49
        pixel_data[50][0] = 4'b0001; // x=0, y=50
        pixel_data[50][1] = 4'b0001; // x=1, y=50
        pixel_data[50][2] = 4'b0001; // x=2, y=50
        pixel_data[50][3] = 4'b0001; // x=3, y=50
        pixel_data[50][4] = 4'b0001; // x=4, y=50
        pixel_data[50][5] = 4'b0001; // x=5, y=50
        pixel_data[50][6] = 4'b0001; // x=6, y=50
        pixel_data[50][7] = 4'b0001; // x=7, y=50
        pixel_data[50][8] = 4'b0001; // x=8, y=50
        pixel_data[50][9] = 4'b0001; // x=9, y=50
        pixel_data[50][10] = 4'b0001; // x=10, y=50
        pixel_data[50][11] = 4'b0001; // x=11, y=50
        pixel_data[50][12] = 4'b0001; // x=12, y=50
        pixel_data[50][13] = 4'b0001; // x=13, y=50
        pixel_data[50][14] = 4'b0001; // x=14, y=50
        pixel_data[50][15] = 4'b0001; // x=15, y=50
        pixel_data[50][16] = 4'b0001; // x=16, y=50
        pixel_data[50][17] = 4'b0001; // x=17, y=50
        pixel_data[50][18] = 4'b0001; // x=18, y=50
        pixel_data[50][19] = 4'b0001; // x=19, y=50
        pixel_data[50][20] = 4'b0001; // x=20, y=50
        pixel_data[50][21] = 4'b0001; // x=21, y=50
        pixel_data[50][22] = 4'b0001; // x=22, y=50
        pixel_data[50][23] = 4'b0001; // x=23, y=50
        pixel_data[50][24] = 4'b0001; // x=24, y=50
        pixel_data[50][25] = 4'b0001; // x=25, y=50
        pixel_data[50][26] = 4'b0001; // x=26, y=50
        pixel_data[50][27] = 4'b0001; // x=27, y=50
        pixel_data[50][28] = 4'b0001; // x=28, y=50
        pixel_data[50][29] = 4'b0001; // x=29, y=50
        pixel_data[50][30] = 4'b0001; // x=30, y=50
        pixel_data[50][31] = 4'b0001; // x=31, y=50
        pixel_data[50][32] = 4'b0001; // x=32, y=50
        pixel_data[50][33] = 4'b0001; // x=33, y=50
        pixel_data[50][34] = 4'b0001; // x=34, y=50
        pixel_data[50][35] = 4'b0001; // x=35, y=50
        pixel_data[50][36] = 4'b0001; // x=36, y=50
        pixel_data[50][37] = 4'b0001; // x=37, y=50
        pixel_data[50][38] = 4'b0001; // x=38, y=50
        pixel_data[50][39] = 4'b0001; // x=39, y=50
        pixel_data[50][40] = 4'b0001; // x=40, y=50
        pixel_data[50][41] = 4'b0001; // x=41, y=50
        pixel_data[50][42] = 4'b0001; // x=42, y=50
        pixel_data[50][43] = 4'b0001; // x=43, y=50
        pixel_data[50][44] = 4'b0001; // x=44, y=50
        pixel_data[50][45] = 4'b0001; // x=45, y=50
        pixel_data[50][46] = 4'b0001; // x=46, y=50
        pixel_data[50][47] = 4'b0001; // x=47, y=50
        pixel_data[50][48] = 4'b0001; // x=48, y=50
        pixel_data[50][49] = 4'b0001; // x=49, y=50
        pixel_data[50][50] = 4'b0001; // x=50, y=50
        pixel_data[50][51] = 4'b0001; // x=51, y=50
        pixel_data[50][52] = 4'b0001; // x=52, y=50
        pixel_data[50][53] = 4'b0001; // x=53, y=50
        pixel_data[50][54] = 4'b0001; // x=54, y=50
        pixel_data[50][55] = 4'b0001; // x=55, y=50
        pixel_data[50][56] = 4'b0001; // x=56, y=50
        pixel_data[50][57] = 4'b0001; // x=57, y=50
        pixel_data[50][58] = 4'b0001; // x=58, y=50
        pixel_data[50][59] = 4'b0001; // x=59, y=50
        pixel_data[51][0] = 4'b0001; // x=0, y=51
        pixel_data[51][1] = 4'b0001; // x=1, y=51
        pixel_data[51][2] = 4'b0001; // x=2, y=51
        pixel_data[51][3] = 4'b0001; // x=3, y=51
        pixel_data[51][4] = 4'b0001; // x=4, y=51
        pixel_data[51][5] = 4'b0001; // x=5, y=51
        pixel_data[51][6] = 4'b0001; // x=6, y=51
        pixel_data[51][7] = 4'b0001; // x=7, y=51
        pixel_data[51][8] = 4'b0001; // x=8, y=51
        pixel_data[51][9] = 4'b0001; // x=9, y=51
        pixel_data[51][10] = 4'b0001; // x=10, y=51
        pixel_data[51][11] = 4'b0001; // x=11, y=51
        pixel_data[51][12] = 4'b0001; // x=12, y=51
        pixel_data[51][13] = 4'b0001; // x=13, y=51
        pixel_data[51][14] = 4'b0001; // x=14, y=51
        pixel_data[51][15] = 4'b0001; // x=15, y=51
        pixel_data[51][16] = 4'b0001; // x=16, y=51
        pixel_data[51][17] = 4'b0001; // x=17, y=51
        pixel_data[51][18] = 4'b0001; // x=18, y=51
        pixel_data[51][19] = 4'b0001; // x=19, y=51
        pixel_data[51][20] = 4'b0001; // x=20, y=51
        pixel_data[51][21] = 4'b0001; // x=21, y=51
        pixel_data[51][22] = 4'b0001; // x=22, y=51
        pixel_data[51][23] = 4'b0001; // x=23, y=51
        pixel_data[51][24] = 4'b0001; // x=24, y=51
        pixel_data[51][25] = 4'b0001; // x=25, y=51
        pixel_data[51][26] = 4'b0001; // x=26, y=51
        pixel_data[51][27] = 4'b0001; // x=27, y=51
        pixel_data[51][28] = 4'b0001; // x=28, y=51
        pixel_data[51][29] = 4'b0001; // x=29, y=51
        pixel_data[51][30] = 4'b0001; // x=30, y=51
        pixel_data[51][31] = 4'b0001; // x=31, y=51
        pixel_data[51][32] = 4'b0001; // x=32, y=51
        pixel_data[51][33] = 4'b0001; // x=33, y=51
        pixel_data[51][34] = 4'b0001; // x=34, y=51
        pixel_data[51][35] = 4'b0001; // x=35, y=51
        pixel_data[51][36] = 4'b0001; // x=36, y=51
        pixel_data[51][37] = 4'b0001; // x=37, y=51
        pixel_data[51][38] = 4'b0001; // x=38, y=51
        pixel_data[51][39] = 4'b0001; // x=39, y=51
        pixel_data[51][40] = 4'b0001; // x=40, y=51
        pixel_data[51][41] = 4'b0001; // x=41, y=51
        pixel_data[51][42] = 4'b0001; // x=42, y=51
        pixel_data[51][43] = 4'b0001; // x=43, y=51
        pixel_data[51][44] = 4'b0001; // x=44, y=51
        pixel_data[51][45] = 4'b0001; // x=45, y=51
        pixel_data[51][46] = 4'b0001; // x=46, y=51
        pixel_data[51][47] = 4'b0001; // x=47, y=51
        pixel_data[51][48] = 4'b0001; // x=48, y=51
        pixel_data[51][49] = 4'b0001; // x=49, y=51
        pixel_data[51][50] = 4'b0001; // x=50, y=51
        pixel_data[51][51] = 4'b0001; // x=51, y=51
        pixel_data[51][52] = 4'b0001; // x=52, y=51
        pixel_data[51][53] = 4'b0001; // x=53, y=51
        pixel_data[51][54] = 4'b0001; // x=54, y=51
        pixel_data[51][55] = 4'b0001; // x=55, y=51
        pixel_data[51][56] = 4'b0001; // x=56, y=51
        pixel_data[51][57] = 4'b0001; // x=57, y=51
        pixel_data[51][58] = 4'b0001; // x=58, y=51
        pixel_data[51][59] = 4'b0001; // x=59, y=51
        pixel_data[52][0] = 4'b0001; // x=0, y=52
        pixel_data[52][1] = 4'b0001; // x=1, y=52
        pixel_data[52][2] = 4'b0001; // x=2, y=52
        pixel_data[52][3] = 4'b0001; // x=3, y=52
        pixel_data[52][4] = 4'b0001; // x=4, y=52
        pixel_data[52][5] = 4'b0001; // x=5, y=52
        pixel_data[52][6] = 4'b0001; // x=6, y=52
        pixel_data[52][7] = 4'b0001; // x=7, y=52
        pixel_data[52][8] = 4'b0001; // x=8, y=52
        pixel_data[52][9] = 4'b0001; // x=9, y=52
        pixel_data[52][10] = 4'b0001; // x=10, y=52
        pixel_data[52][11] = 4'b0001; // x=11, y=52
        pixel_data[52][12] = 4'b0001; // x=12, y=52
        pixel_data[52][13] = 4'b0001; // x=13, y=52
        pixel_data[52][14] = 4'b0001; // x=14, y=52
        pixel_data[52][15] = 4'b0001; // x=15, y=52
        pixel_data[52][16] = 4'b0001; // x=16, y=52
        pixel_data[52][17] = 4'b0001; // x=17, y=52
        pixel_data[52][18] = 4'b0001; // x=18, y=52
        pixel_data[52][19] = 4'b0001; // x=19, y=52
        pixel_data[52][20] = 4'b0001; // x=20, y=52
        pixel_data[52][21] = 4'b0001; // x=21, y=52
        pixel_data[52][22] = 4'b0001; // x=22, y=52
        pixel_data[52][23] = 4'b0001; // x=23, y=52
        pixel_data[52][24] = 4'b0001; // x=24, y=52
        pixel_data[52][25] = 4'b0001; // x=25, y=52
        pixel_data[52][26] = 4'b0001; // x=26, y=52
        pixel_data[52][27] = 4'b0001; // x=27, y=52
        pixel_data[52][28] = 4'b0001; // x=28, y=52
        pixel_data[52][29] = 4'b0001; // x=29, y=52
        pixel_data[52][30] = 4'b0001; // x=30, y=52
        pixel_data[52][31] = 4'b0001; // x=31, y=52
        pixel_data[52][32] = 4'b0001; // x=32, y=52
        pixel_data[52][33] = 4'b0001; // x=33, y=52
        pixel_data[52][34] = 4'b0001; // x=34, y=52
        pixel_data[52][35] = 4'b0001; // x=35, y=52
        pixel_data[52][36] = 4'b0001; // x=36, y=52
        pixel_data[52][37] = 4'b0001; // x=37, y=52
        pixel_data[52][38] = 4'b0001; // x=38, y=52
        pixel_data[52][39] = 4'b0001; // x=39, y=52
        pixel_data[52][40] = 4'b0001; // x=40, y=52
        pixel_data[52][41] = 4'b0001; // x=41, y=52
        pixel_data[52][42] = 4'b0001; // x=42, y=52
        pixel_data[52][43] = 4'b0001; // x=43, y=52
        pixel_data[52][44] = 4'b0001; // x=44, y=52
        pixel_data[52][45] = 4'b0001; // x=45, y=52
        pixel_data[52][46] = 4'b0001; // x=46, y=52
        pixel_data[52][47] = 4'b0001; // x=47, y=52
        pixel_data[52][48] = 4'b0001; // x=48, y=52
        pixel_data[52][49] = 4'b0001; // x=49, y=52
        pixel_data[52][50] = 4'b0001; // x=50, y=52
        pixel_data[52][51] = 4'b0001; // x=51, y=52
        pixel_data[52][52] = 4'b0001; // x=52, y=52
        pixel_data[52][53] = 4'b0001; // x=53, y=52
        pixel_data[52][54] = 4'b0001; // x=54, y=52
        pixel_data[52][55] = 4'b0001; // x=55, y=52
        pixel_data[52][56] = 4'b0001; // x=56, y=52
        pixel_data[52][57] = 4'b0001; // x=57, y=52
        pixel_data[52][58] = 4'b0001; // x=58, y=52
        pixel_data[52][59] = 4'b0001; // x=59, y=52
        pixel_data[53][0] = 4'b0001; // x=0, y=53
        pixel_data[53][1] = 4'b0001; // x=1, y=53
        pixel_data[53][2] = 4'b0001; // x=2, y=53
        pixel_data[53][3] = 4'b0001; // x=3, y=53
        pixel_data[53][4] = 4'b0001; // x=4, y=53
        pixel_data[53][5] = 4'b0001; // x=5, y=53
        pixel_data[53][6] = 4'b0001; // x=6, y=53
        pixel_data[53][7] = 4'b0001; // x=7, y=53
        pixel_data[53][8] = 4'b0001; // x=8, y=53
        pixel_data[53][9] = 4'b0001; // x=9, y=53
        pixel_data[53][10] = 4'b0001; // x=10, y=53
        pixel_data[53][11] = 4'b0001; // x=11, y=53
        pixel_data[53][12] = 4'b0001; // x=12, y=53
        pixel_data[53][13] = 4'b0001; // x=13, y=53
        pixel_data[53][14] = 4'b0001; // x=14, y=53
        pixel_data[53][15] = 4'b0001; // x=15, y=53
        pixel_data[53][16] = 4'b0001; // x=16, y=53
        pixel_data[53][17] = 4'b0001; // x=17, y=53
        pixel_data[53][18] = 4'b0001; // x=18, y=53
        pixel_data[53][19] = 4'b0001; // x=19, y=53
        pixel_data[53][20] = 4'b0001; // x=20, y=53
        pixel_data[53][21] = 4'b0001; // x=21, y=53
        pixel_data[53][22] = 4'b0001; // x=22, y=53
        pixel_data[53][23] = 4'b0001; // x=23, y=53
        pixel_data[53][24] = 4'b0001; // x=24, y=53
        pixel_data[53][25] = 4'b0001; // x=25, y=53
        pixel_data[53][26] = 4'b0001; // x=26, y=53
        pixel_data[53][27] = 4'b0001; // x=27, y=53
        pixel_data[53][28] = 4'b0001; // x=28, y=53
        pixel_data[53][29] = 4'b0001; // x=29, y=53
        pixel_data[53][30] = 4'b0001; // x=30, y=53
        pixel_data[53][31] = 4'b0001; // x=31, y=53
        pixel_data[53][32] = 4'b0001; // x=32, y=53
        pixel_data[53][33] = 4'b0001; // x=33, y=53
        pixel_data[53][34] = 4'b0001; // x=34, y=53
        pixel_data[53][35] = 4'b0001; // x=35, y=53
        pixel_data[53][36] = 4'b0001; // x=36, y=53
        pixel_data[53][37] = 4'b0001; // x=37, y=53
        pixel_data[53][38] = 4'b0001; // x=38, y=53
        pixel_data[53][39] = 4'b0001; // x=39, y=53
        pixel_data[53][40] = 4'b0001; // x=40, y=53
        pixel_data[53][41] = 4'b0001; // x=41, y=53
        pixel_data[53][42] = 4'b0001; // x=42, y=53
        pixel_data[53][43] = 4'b0001; // x=43, y=53
        pixel_data[53][44] = 4'b0001; // x=44, y=53
        pixel_data[53][45] = 4'b0001; // x=45, y=53
        pixel_data[53][46] = 4'b0001; // x=46, y=53
        pixel_data[53][47] = 4'b0001; // x=47, y=53
        pixel_data[53][48] = 4'b0001; // x=48, y=53
        pixel_data[53][49] = 4'b0001; // x=49, y=53
        pixel_data[53][50] = 4'b0001; // x=50, y=53
        pixel_data[53][51] = 4'b0001; // x=51, y=53
        pixel_data[53][52] = 4'b0001; // x=52, y=53
        pixel_data[53][53] = 4'b0001; // x=53, y=53
        pixel_data[53][54] = 4'b0001; // x=54, y=53
        pixel_data[53][55] = 4'b0001; // x=55, y=53
        pixel_data[53][56] = 4'b0001; // x=56, y=53
        pixel_data[53][57] = 4'b0001; // x=57, y=53
        pixel_data[53][58] = 4'b0001; // x=58, y=53
        pixel_data[53][59] = 4'b0001; // x=59, y=53
        pixel_data[54][0] = 4'b0001; // x=0, y=54
        pixel_data[54][1] = 4'b0001; // x=1, y=54
        pixel_data[54][2] = 4'b0001; // x=2, y=54
        pixel_data[54][3] = 4'b0001; // x=3, y=54
        pixel_data[54][4] = 4'b0001; // x=4, y=54
        pixel_data[54][5] = 4'b0001; // x=5, y=54
        pixel_data[54][6] = 4'b0001; // x=6, y=54
        pixel_data[54][7] = 4'b0001; // x=7, y=54
        pixel_data[54][8] = 4'b0001; // x=8, y=54
        pixel_data[54][9] = 4'b0001; // x=9, y=54
        pixel_data[54][10] = 4'b0001; // x=10, y=54
        pixel_data[54][11] = 4'b0001; // x=11, y=54
        pixel_data[54][12] = 4'b0001; // x=12, y=54
        pixel_data[54][13] = 4'b0001; // x=13, y=54
        pixel_data[54][14] = 4'b0001; // x=14, y=54
        pixel_data[54][15] = 4'b0001; // x=15, y=54
        pixel_data[54][16] = 4'b0001; // x=16, y=54
        pixel_data[54][17] = 4'b0001; // x=17, y=54
        pixel_data[54][18] = 4'b0001; // x=18, y=54
        pixel_data[54][19] = 4'b0001; // x=19, y=54
        pixel_data[54][20] = 4'b0001; // x=20, y=54
        pixel_data[54][21] = 4'b0001; // x=21, y=54
        pixel_data[54][22] = 4'b0001; // x=22, y=54
        pixel_data[54][23] = 4'b0001; // x=23, y=54
        pixel_data[54][24] = 4'b0001; // x=24, y=54
        pixel_data[54][25] = 4'b0001; // x=25, y=54
        pixel_data[54][26] = 4'b0001; // x=26, y=54
        pixel_data[54][27] = 4'b0001; // x=27, y=54
        pixel_data[54][28] = 4'b0001; // x=28, y=54
        pixel_data[54][29] = 4'b0001; // x=29, y=54
        pixel_data[54][30] = 4'b0001; // x=30, y=54
        pixel_data[54][31] = 4'b0001; // x=31, y=54
        pixel_data[54][32] = 4'b0001; // x=32, y=54
        pixel_data[54][33] = 4'b0001; // x=33, y=54
        pixel_data[54][34] = 4'b0001; // x=34, y=54
        pixel_data[54][35] = 4'b0001; // x=35, y=54
        pixel_data[54][36] = 4'b0001; // x=36, y=54
        pixel_data[54][37] = 4'b0001; // x=37, y=54
        pixel_data[54][38] = 4'b0001; // x=38, y=54
        pixel_data[54][39] = 4'b0001; // x=39, y=54
        pixel_data[54][40] = 4'b0001; // x=40, y=54
        pixel_data[54][41] = 4'b0001; // x=41, y=54
        pixel_data[54][42] = 4'b0001; // x=42, y=54
        pixel_data[54][43] = 4'b0001; // x=43, y=54
        pixel_data[54][44] = 4'b0001; // x=44, y=54
        pixel_data[54][45] = 4'b0001; // x=45, y=54
        pixel_data[54][46] = 4'b0001; // x=46, y=54
        pixel_data[54][47] = 4'b0001; // x=47, y=54
        pixel_data[54][48] = 4'b0001; // x=48, y=54
        pixel_data[54][49] = 4'b0001; // x=49, y=54
        pixel_data[54][50] = 4'b0001; // x=50, y=54
        pixel_data[54][51] = 4'b0001; // x=51, y=54
        pixel_data[54][52] = 4'b0001; // x=52, y=54
        pixel_data[54][53] = 4'b0001; // x=53, y=54
        pixel_data[54][54] = 4'b0001; // x=54, y=54
        pixel_data[54][55] = 4'b0001; // x=55, y=54
        pixel_data[54][56] = 4'b0001; // x=56, y=54
        pixel_data[54][57] = 4'b0001; // x=57, y=54
        pixel_data[54][58] = 4'b0001; // x=58, y=54
        pixel_data[54][59] = 4'b0001; // x=59, y=54
        pixel_data[55][0] = 4'b0001; // x=0, y=55
        pixel_data[55][1] = 4'b0001; // x=1, y=55
        pixel_data[55][2] = 4'b0001; // x=2, y=55
        pixel_data[55][3] = 4'b0001; // x=3, y=55
        pixel_data[55][4] = 4'b0001; // x=4, y=55
        pixel_data[55][5] = 4'b0001; // x=5, y=55
        pixel_data[55][6] = 4'b0001; // x=6, y=55
        pixel_data[55][7] = 4'b0001; // x=7, y=55
        pixel_data[55][8] = 4'b0001; // x=8, y=55
        pixel_data[55][9] = 4'b0001; // x=9, y=55
        pixel_data[55][10] = 4'b0001; // x=10, y=55
        pixel_data[55][11] = 4'b0001; // x=11, y=55
        pixel_data[55][12] = 4'b0001; // x=12, y=55
        pixel_data[55][13] = 4'b0001; // x=13, y=55
        pixel_data[55][14] = 4'b0001; // x=14, y=55
        pixel_data[55][15] = 4'b0001; // x=15, y=55
        pixel_data[55][16] = 4'b0001; // x=16, y=55
        pixel_data[55][17] = 4'b0001; // x=17, y=55
        pixel_data[55][18] = 4'b0001; // x=18, y=55
        pixel_data[55][19] = 4'b0001; // x=19, y=55
        pixel_data[55][20] = 4'b0001; // x=20, y=55
        pixel_data[55][21] = 4'b0001; // x=21, y=55
        pixel_data[55][22] = 4'b0001; // x=22, y=55
        pixel_data[55][23] = 4'b0001; // x=23, y=55
        pixel_data[55][24] = 4'b0001; // x=24, y=55
        pixel_data[55][25] = 4'b0001; // x=25, y=55
        pixel_data[55][26] = 4'b0001; // x=26, y=55
        pixel_data[55][27] = 4'b0001; // x=27, y=55
        pixel_data[55][28] = 4'b0001; // x=28, y=55
        pixel_data[55][29] = 4'b0001; // x=29, y=55
        pixel_data[55][30] = 4'b0001; // x=30, y=55
        pixel_data[55][31] = 4'b0001; // x=31, y=55
        pixel_data[55][32] = 4'b0001; // x=32, y=55
        pixel_data[55][33] = 4'b0001; // x=33, y=55
        pixel_data[55][34] = 4'b0001; // x=34, y=55
        pixel_data[55][35] = 4'b0001; // x=35, y=55
        pixel_data[55][36] = 4'b0001; // x=36, y=55
        pixel_data[55][37] = 4'b0001; // x=37, y=55
        pixel_data[55][38] = 4'b0001; // x=38, y=55
        pixel_data[55][39] = 4'b0001; // x=39, y=55
        pixel_data[55][40] = 4'b0001; // x=40, y=55
        pixel_data[55][41] = 4'b0001; // x=41, y=55
        pixel_data[55][42] = 4'b0001; // x=42, y=55
        pixel_data[55][43] = 4'b0001; // x=43, y=55
        pixel_data[55][44] = 4'b0001; // x=44, y=55
        pixel_data[55][45] = 4'b0001; // x=45, y=55
        pixel_data[55][46] = 4'b0001; // x=46, y=55
        pixel_data[55][47] = 4'b0001; // x=47, y=55
        pixel_data[55][48] = 4'b0001; // x=48, y=55
        pixel_data[55][49] = 4'b0001; // x=49, y=55
        pixel_data[55][50] = 4'b0001; // x=50, y=55
        pixel_data[55][51] = 4'b0001; // x=51, y=55
        pixel_data[55][52] = 4'b0001; // x=52, y=55
        pixel_data[55][53] = 4'b0001; // x=53, y=55
        pixel_data[55][54] = 4'b0001; // x=54, y=55
        pixel_data[55][55] = 4'b0001; // x=55, y=55
        pixel_data[55][56] = 4'b0001; // x=56, y=55
        pixel_data[55][57] = 4'b0001; // x=57, y=55
        pixel_data[55][58] = 4'b0001; // x=58, y=55
        pixel_data[55][59] = 4'b0001; // x=59, y=55
        pixel_data[56][0] = 4'b0001; // x=0, y=56
        pixel_data[56][1] = 4'b0001; // x=1, y=56
        pixel_data[56][2] = 4'b0001; // x=2, y=56
        pixel_data[56][3] = 4'b0001; // x=3, y=56
        pixel_data[56][4] = 4'b0001; // x=4, y=56
        pixel_data[56][5] = 4'b0001; // x=5, y=56
        pixel_data[56][6] = 4'b0001; // x=6, y=56
        pixel_data[56][7] = 4'b0001; // x=7, y=56
        pixel_data[56][8] = 4'b0001; // x=8, y=56
        pixel_data[56][9] = 4'b0001; // x=9, y=56
        pixel_data[56][10] = 4'b0001; // x=10, y=56
        pixel_data[56][11] = 4'b0001; // x=11, y=56
        pixel_data[56][12] = 4'b0001; // x=12, y=56
        pixel_data[56][13] = 4'b0001; // x=13, y=56
        pixel_data[56][14] = 4'b0001; // x=14, y=56
        pixel_data[56][15] = 4'b0001; // x=15, y=56
        pixel_data[56][16] = 4'b0001; // x=16, y=56
        pixel_data[56][17] = 4'b0001; // x=17, y=56
        pixel_data[56][18] = 4'b0001; // x=18, y=56
        pixel_data[56][19] = 4'b0001; // x=19, y=56
        pixel_data[56][20] = 4'b0001; // x=20, y=56
        pixel_data[56][21] = 4'b0001; // x=21, y=56
        pixel_data[56][22] = 4'b0001; // x=22, y=56
        pixel_data[56][23] = 4'b0001; // x=23, y=56
        pixel_data[56][24] = 4'b0001; // x=24, y=56
        pixel_data[56][25] = 4'b0001; // x=25, y=56
        pixel_data[56][26] = 4'b0001; // x=26, y=56
        pixel_data[56][27] = 4'b0001; // x=27, y=56
        pixel_data[56][28] = 4'b0001; // x=28, y=56
        pixel_data[56][29] = 4'b0001; // x=29, y=56
        pixel_data[56][30] = 4'b0001; // x=30, y=56
        pixel_data[56][31] = 4'b0001; // x=31, y=56
        pixel_data[56][32] = 4'b0001; // x=32, y=56
        pixel_data[56][33] = 4'b0001; // x=33, y=56
        pixel_data[56][34] = 4'b0001; // x=34, y=56
        pixel_data[56][35] = 4'b0001; // x=35, y=56
        pixel_data[56][36] = 4'b0001; // x=36, y=56
        pixel_data[56][37] = 4'b0001; // x=37, y=56
        pixel_data[56][38] = 4'b0001; // x=38, y=56
        pixel_data[56][39] = 4'b0001; // x=39, y=56
        pixel_data[56][40] = 4'b0001; // x=40, y=56
        pixel_data[56][41] = 4'b0001; // x=41, y=56
        pixel_data[56][42] = 4'b0001; // x=42, y=56
        pixel_data[56][43] = 4'b0001; // x=43, y=56
        pixel_data[56][44] = 4'b0001; // x=44, y=56
        pixel_data[56][45] = 4'b0001; // x=45, y=56
        pixel_data[56][46] = 4'b0001; // x=46, y=56
        pixel_data[56][47] = 4'b0001; // x=47, y=56
        pixel_data[56][48] = 4'b0001; // x=48, y=56
        pixel_data[56][49] = 4'b0001; // x=49, y=56
        pixel_data[56][50] = 4'b0001; // x=50, y=56
        pixel_data[56][51] = 4'b0001; // x=51, y=56
        pixel_data[56][52] = 4'b0001; // x=52, y=56
        pixel_data[56][53] = 4'b0001; // x=53, y=56
        pixel_data[56][54] = 4'b0001; // x=54, y=56
        pixel_data[56][55] = 4'b0001; // x=55, y=56
        pixel_data[56][56] = 4'b0001; // x=56, y=56
        pixel_data[56][57] = 4'b0001; // x=57, y=56
        pixel_data[56][58] = 4'b0001; // x=58, y=56
        pixel_data[56][59] = 4'b0001; // x=59, y=56
        pixel_data[57][0] = 4'b0001; // x=0, y=57
        pixel_data[57][1] = 4'b0001; // x=1, y=57
        pixel_data[57][2] = 4'b0001; // x=2, y=57
        pixel_data[57][3] = 4'b0001; // x=3, y=57
        pixel_data[57][4] = 4'b0001; // x=4, y=57
        pixel_data[57][5] = 4'b0001; // x=5, y=57
        pixel_data[57][6] = 4'b0001; // x=6, y=57
        pixel_data[57][7] = 4'b0001; // x=7, y=57
        pixel_data[57][8] = 4'b0001; // x=8, y=57
        pixel_data[57][9] = 4'b0001; // x=9, y=57
        pixel_data[57][10] = 4'b0001; // x=10, y=57
        pixel_data[57][11] = 4'b0001; // x=11, y=57
        pixel_data[57][12] = 4'b0001; // x=12, y=57
        pixel_data[57][13] = 4'b0001; // x=13, y=57
        pixel_data[57][14] = 4'b0001; // x=14, y=57
        pixel_data[57][15] = 4'b0001; // x=15, y=57
        pixel_data[57][16] = 4'b0001; // x=16, y=57
        pixel_data[57][17] = 4'b0001; // x=17, y=57
        pixel_data[57][18] = 4'b0001; // x=18, y=57
        pixel_data[57][19] = 4'b0001; // x=19, y=57
        pixel_data[57][20] = 4'b0001; // x=20, y=57
        pixel_data[57][21] = 4'b0001; // x=21, y=57
        pixel_data[57][22] = 4'b0001; // x=22, y=57
        pixel_data[57][23] = 4'b0001; // x=23, y=57
        pixel_data[57][24] = 4'b0001; // x=24, y=57
        pixel_data[57][25] = 4'b0001; // x=25, y=57
        pixel_data[57][26] = 4'b0001; // x=26, y=57
        pixel_data[57][27] = 4'b0001; // x=27, y=57
        pixel_data[57][28] = 4'b0001; // x=28, y=57
        pixel_data[57][29] = 4'b0001; // x=29, y=57
        pixel_data[57][30] = 4'b0001; // x=30, y=57
        pixel_data[57][31] = 4'b0001; // x=31, y=57
        pixel_data[57][32] = 4'b0001; // x=32, y=57
        pixel_data[57][33] = 4'b0001; // x=33, y=57
        pixel_data[57][34] = 4'b0001; // x=34, y=57
        pixel_data[57][35] = 4'b0001; // x=35, y=57
        pixel_data[57][36] = 4'b0001; // x=36, y=57
        pixel_data[57][37] = 4'b0001; // x=37, y=57
        pixel_data[57][38] = 4'b0001; // x=38, y=57
        pixel_data[57][39] = 4'b0001; // x=39, y=57
        pixel_data[57][40] = 4'b0001; // x=40, y=57
        pixel_data[57][41] = 4'b0001; // x=41, y=57
        pixel_data[57][42] = 4'b0001; // x=42, y=57
        pixel_data[57][43] = 4'b0001; // x=43, y=57
        pixel_data[57][44] = 4'b0001; // x=44, y=57
        pixel_data[57][45] = 4'b0001; // x=45, y=57
        pixel_data[57][46] = 4'b0001; // x=46, y=57
        pixel_data[57][47] = 4'b0001; // x=47, y=57
        pixel_data[57][48] = 4'b0001; // x=48, y=57
        pixel_data[57][49] = 4'b0001; // x=49, y=57
        pixel_data[57][50] = 4'b0001; // x=50, y=57
        pixel_data[57][51] = 4'b0001; // x=51, y=57
        pixel_data[57][52] = 4'b0001; // x=52, y=57
        pixel_data[57][53] = 4'b0001; // x=53, y=57
        pixel_data[57][54] = 4'b0001; // x=54, y=57
        pixel_data[57][55] = 4'b0001; // x=55, y=57
        pixel_data[57][56] = 4'b0001; // x=56, y=57
        pixel_data[57][57] = 4'b0001; // x=57, y=57
        pixel_data[57][58] = 4'b0001; // x=58, y=57
        pixel_data[57][59] = 4'b0001; // x=59, y=57
        pixel_data[58][0] = 4'b0001; // x=0, y=58
        pixel_data[58][1] = 4'b0001; // x=1, y=58
        pixel_data[58][2] = 4'b0001; // x=2, y=58
        pixel_data[58][3] = 4'b0001; // x=3, y=58
        pixel_data[58][4] = 4'b0001; // x=4, y=58
        pixel_data[58][5] = 4'b0001; // x=5, y=58
        pixel_data[58][6] = 4'b0001; // x=6, y=58
        pixel_data[58][7] = 4'b0001; // x=7, y=58
        pixel_data[58][8] = 4'b0001; // x=8, y=58
        pixel_data[58][9] = 4'b0001; // x=9, y=58
        pixel_data[58][10] = 4'b0001; // x=10, y=58
        pixel_data[58][11] = 4'b0001; // x=11, y=58
        pixel_data[58][12] = 4'b0001; // x=12, y=58
        pixel_data[58][13] = 4'b0001; // x=13, y=58
        pixel_data[58][14] = 4'b0001; // x=14, y=58
        pixel_data[58][15] = 4'b0001; // x=15, y=58
        pixel_data[58][16] = 4'b0001; // x=16, y=58
        pixel_data[58][17] = 4'b0001; // x=17, y=58
        pixel_data[58][18] = 4'b0001; // x=18, y=58
        pixel_data[58][19] = 4'b0001; // x=19, y=58
        pixel_data[58][20] = 4'b0001; // x=20, y=58
        pixel_data[58][21] = 4'b0001; // x=21, y=58
        pixel_data[58][22] = 4'b0001; // x=22, y=58
        pixel_data[58][23] = 4'b0001; // x=23, y=58
        pixel_data[58][24] = 4'b0001; // x=24, y=58
        pixel_data[58][25] = 4'b0001; // x=25, y=58
        pixel_data[58][26] = 4'b0001; // x=26, y=58
        pixel_data[58][27] = 4'b0001; // x=27, y=58
        pixel_data[58][28] = 4'b0001; // x=28, y=58
        pixel_data[58][29] = 4'b0001; // x=29, y=58
        pixel_data[58][30] = 4'b0001; // x=30, y=58
        pixel_data[58][31] = 4'b0001; // x=31, y=58
        pixel_data[58][32] = 4'b0001; // x=32, y=58
        pixel_data[58][33] = 4'b0001; // x=33, y=58
        pixel_data[58][34] = 4'b0001; // x=34, y=58
        pixel_data[58][35] = 4'b0001; // x=35, y=58
        pixel_data[58][36] = 4'b0001; // x=36, y=58
        pixel_data[58][37] = 4'b0001; // x=37, y=58
        pixel_data[58][38] = 4'b0001; // x=38, y=58
        pixel_data[58][39] = 4'b0001; // x=39, y=58
        pixel_data[58][40] = 4'b0001; // x=40, y=58
        pixel_data[58][41] = 4'b0001; // x=41, y=58
        pixel_data[58][42] = 4'b0001; // x=42, y=58
        pixel_data[58][43] = 4'b0001; // x=43, y=58
        pixel_data[58][44] = 4'b0001; // x=44, y=58
        pixel_data[58][45] = 4'b0001; // x=45, y=58
        pixel_data[58][46] = 4'b0001; // x=46, y=58
        pixel_data[58][47] = 4'b0001; // x=47, y=58
        pixel_data[58][48] = 4'b0001; // x=48, y=58
        pixel_data[58][49] = 4'b0001; // x=49, y=58
        pixel_data[58][50] = 4'b0001; // x=50, y=58
        pixel_data[58][51] = 4'b0001; // x=51, y=58
        pixel_data[58][52] = 4'b0001; // x=52, y=58
        pixel_data[58][53] = 4'b0001; // x=53, y=58
        pixel_data[58][54] = 4'b0001; // x=54, y=58
        pixel_data[58][55] = 4'b0001; // x=55, y=58
        pixel_data[58][56] = 4'b0001; // x=56, y=58
        pixel_data[58][57] = 4'b0001; // x=57, y=58
        pixel_data[58][58] = 4'b0001; // x=58, y=58
        pixel_data[58][59] = 4'b0001; // x=59, y=58
        pixel_data[59][0] = 4'b0001; // x=0, y=59
        pixel_data[59][1] = 4'b0001; // x=1, y=59
        pixel_data[59][2] = 4'b0001; // x=2, y=59
        pixel_data[59][3] = 4'b0001; // x=3, y=59
        pixel_data[59][4] = 4'b0001; // x=4, y=59
        pixel_data[59][5] = 4'b0001; // x=5, y=59
        pixel_data[59][6] = 4'b0001; // x=6, y=59
        pixel_data[59][7] = 4'b0001; // x=7, y=59
        pixel_data[59][8] = 4'b0001; // x=8, y=59
        pixel_data[59][9] = 4'b0001; // x=9, y=59
        pixel_data[59][10] = 4'b0001; // x=10, y=59
        pixel_data[59][11] = 4'b0001; // x=11, y=59
        pixel_data[59][12] = 4'b0001; // x=12, y=59
        pixel_data[59][13] = 4'b0001; // x=13, y=59
        pixel_data[59][14] = 4'b0001; // x=14, y=59
        pixel_data[59][15] = 4'b0001; // x=15, y=59
        pixel_data[59][16] = 4'b0001; // x=16, y=59
        pixel_data[59][17] = 4'b0001; // x=17, y=59
        pixel_data[59][18] = 4'b0001; // x=18, y=59
        pixel_data[59][19] = 4'b0001; // x=19, y=59
        pixel_data[59][20] = 4'b0001; // x=20, y=59
        pixel_data[59][21] = 4'b0001; // x=21, y=59
        pixel_data[59][22] = 4'b0001; // x=22, y=59
        pixel_data[59][23] = 4'b0001; // x=23, y=59
        pixel_data[59][24] = 4'b0001; // x=24, y=59
        pixel_data[59][25] = 4'b0001; // x=25, y=59
        pixel_data[59][26] = 4'b0001; // x=26, y=59
        pixel_data[59][27] = 4'b0001; // x=27, y=59
        pixel_data[59][28] = 4'b0001; // x=28, y=59
        pixel_data[59][29] = 4'b0001; // x=29, y=59
        pixel_data[59][30] = 4'b0001; // x=30, y=59
        pixel_data[59][31] = 4'b0001; // x=31, y=59
        pixel_data[59][32] = 4'b0001; // x=32, y=59
        pixel_data[59][33] = 4'b0001; // x=33, y=59
        pixel_data[59][34] = 4'b0001; // x=34, y=59
        pixel_data[59][35] = 4'b0001; // x=35, y=59
        pixel_data[59][36] = 4'b0001; // x=36, y=59
        pixel_data[59][37] = 4'b0001; // x=37, y=59
        pixel_data[59][38] = 4'b0001; // x=38, y=59
        pixel_data[59][39] = 4'b0001; // x=39, y=59
        pixel_data[59][40] = 4'b0001; // x=40, y=59
        pixel_data[59][41] = 4'b0001; // x=41, y=59
        pixel_data[59][42] = 4'b0001; // x=42, y=59
        pixel_data[59][43] = 4'b0001; // x=43, y=59
        pixel_data[59][44] = 4'b0001; // x=44, y=59
        pixel_data[59][45] = 4'b0001; // x=45, y=59
        pixel_data[59][46] = 4'b0001; // x=46, y=59
        pixel_data[59][47] = 4'b0001; // x=47, y=59
        pixel_data[59][48] = 4'b0001; // x=48, y=59
        pixel_data[59][49] = 4'b0001; // x=49, y=59
        pixel_data[59][50] = 4'b0001; // x=50, y=59
        pixel_data[59][51] = 4'b0001; // x=51, y=59
        pixel_data[59][52] = 4'b0001; // x=52, y=59
        pixel_data[59][53] = 4'b0001; // x=53, y=59
        pixel_data[59][54] = 4'b0001; // x=54, y=59
        pixel_data[59][55] = 4'b0001; // x=55, y=59
        pixel_data[59][56] = 4'b0001; // x=56, y=59
        pixel_data[59][57] = 4'b0001; // x=57, y=59
        pixel_data[59][58] = 4'b0001; // x=58, y=59
        pixel_data[59][59] = 4'b0001; // x=59, y=59
    end
endmodule

